magic
tech sky130A
magscale 1 2
timestamp 1633951243
<< locali >>
rect 3617 16507 3651 16745
rect 6745 13787 6779 13957
rect 16589 13175 16623 13345
rect 12449 9503 12483 9673
rect 19901 5083 19935 5253
rect 21557 3655 21591 14229
rect 21649 3927 21683 4981
rect 12817 3383 12851 3485
rect 16497 2907 16531 3077
rect 16681 2839 16715 3009
<< viali >>
rect 6377 22117 6411 22151
rect 4169 22049 4203 22083
rect 6837 22049 6871 22083
rect 7941 22049 7975 22083
rect 11529 22049 11563 22083
rect 14841 22049 14875 22083
rect 17325 22049 17359 22083
rect 19901 22049 19935 22083
rect 1869 21981 1903 22015
rect 3065 21981 3099 22015
rect 4445 21981 4479 22015
rect 5641 21981 5675 22015
rect 6561 21981 6595 22015
rect 6653 21981 6687 22015
rect 6929 21981 6963 22015
rect 7757 21981 7791 22015
rect 9413 21981 9447 22015
rect 10057 21981 10091 22015
rect 10793 21981 10827 22015
rect 10977 21981 11011 22015
rect 11805 21981 11839 22015
rect 12909 21981 12943 22015
rect 14197 21981 14231 22015
rect 15117 21981 15151 22015
rect 17141 21981 17175 22015
rect 18521 21981 18555 22015
rect 19441 21981 19475 22015
rect 20177 21981 20211 22015
rect 3249 21913 3283 21947
rect 14381 21913 14415 21947
rect 1961 21845 1995 21879
rect 5733 21845 5767 21879
rect 9505 21845 9539 21879
rect 10241 21845 10275 21879
rect 10885 21845 10919 21879
rect 13001 21845 13035 21879
rect 18613 21845 18647 21879
rect 19257 21845 19291 21879
rect 4261 21641 4295 21675
rect 4997 21641 5031 21675
rect 5181 21641 5215 21675
rect 6745 21641 6779 21675
rect 8401 21641 8435 21675
rect 9505 21641 9539 21675
rect 11713 21641 11747 21675
rect 12449 21641 12483 21675
rect 17877 21641 17911 21675
rect 1869 21573 1903 21607
rect 2053 21573 2087 21607
rect 6837 21573 6871 21607
rect 13369 21573 13403 21607
rect 15945 21573 15979 21607
rect 16865 21573 16899 21607
rect 18613 21573 18647 21607
rect 2513 21505 2547 21539
rect 4169 21505 4203 21539
rect 5178 21505 5212 21539
rect 5641 21505 5675 21539
rect 6561 21505 6595 21539
rect 8309 21505 8343 21539
rect 9413 21505 9447 21539
rect 10241 21505 10275 21539
rect 11621 21505 11655 21539
rect 12265 21505 12299 21539
rect 12541 21505 12575 21539
rect 14197 21505 14231 21539
rect 14381 21505 14415 21539
rect 14841 21505 14875 21539
rect 15025 21505 15059 21539
rect 15117 21505 15151 21539
rect 15209 21505 15243 21539
rect 17693 21505 17727 21539
rect 17969 21505 18003 21539
rect 18429 21505 18463 21539
rect 19257 21505 19291 21539
rect 19901 21505 19935 21539
rect 4445 21437 4479 21471
rect 5549 21437 5583 21471
rect 6377 21437 6411 21471
rect 6929 21437 6963 21471
rect 8493 21437 8527 21471
rect 10517 21437 10551 21471
rect 13461 21437 13495 21471
rect 13553 21437 13587 21471
rect 16129 21437 16163 21471
rect 20177 21437 20211 21471
rect 2697 21369 2731 21403
rect 7941 21369 7975 21403
rect 13001 21369 13035 21403
rect 17049 21369 17083 21403
rect 19349 21369 19383 21403
rect 3801 21301 3835 21335
rect 10057 21301 10091 21335
rect 10425 21301 10459 21335
rect 12265 21301 12299 21335
rect 14197 21301 14231 21335
rect 15393 21301 15427 21335
rect 17509 21301 17543 21335
rect 18797 21301 18831 21335
rect 1961 21097 1995 21131
rect 6929 21097 6963 21131
rect 7941 21097 7975 21131
rect 9321 21097 9355 21131
rect 11713 21097 11747 21131
rect 12909 21097 12943 21131
rect 13461 21097 13495 21131
rect 14381 21097 14415 21131
rect 16405 21097 16439 21131
rect 2789 21029 2823 21063
rect 3801 21029 3835 21063
rect 7849 21029 7883 21063
rect 9965 21029 9999 21063
rect 11897 21029 11931 21063
rect 17325 21029 17359 21063
rect 4353 20961 4387 20995
rect 9505 20961 9539 20995
rect 10609 20961 10643 20995
rect 11805 20961 11839 20995
rect 15025 20961 15059 20995
rect 16497 20961 16531 20995
rect 16589 20961 16623 20995
rect 17785 20961 17819 20995
rect 17877 20961 17911 20995
rect 5273 20893 5307 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6009 20893 6043 20927
rect 6147 20893 6181 20927
rect 6837 20893 6871 20927
rect 7757 20893 7791 20927
rect 8033 20893 8067 20927
rect 8217 20893 8251 20927
rect 9229 20893 9263 20927
rect 10333 20893 10367 20927
rect 12173 20893 12207 20927
rect 13090 20893 13124 20927
rect 13553 20893 13587 20927
rect 16681 20893 16715 20927
rect 16865 20893 16899 20927
rect 18521 20893 18555 20927
rect 19625 20893 19659 20927
rect 20453 20893 20487 20927
rect 1869 20825 1903 20859
rect 2605 20825 2639 20859
rect 5089 20825 5123 20859
rect 9505 20825 9539 20859
rect 14749 20825 14783 20859
rect 18613 20825 18647 20859
rect 4169 20757 4203 20791
rect 4261 20757 4295 20791
rect 6285 20757 6319 20791
rect 7481 20757 7515 20791
rect 10425 20757 10459 20791
rect 11437 20757 11471 20791
rect 12081 20757 12115 20791
rect 13093 20757 13127 20791
rect 14841 20757 14875 20791
rect 16129 20757 16163 20791
rect 17693 20757 17727 20791
rect 19809 20757 19843 20791
rect 20637 20757 20671 20791
rect 2329 20553 2363 20587
rect 3709 20553 3743 20587
rect 8677 20553 8711 20587
rect 10977 20553 11011 20587
rect 11621 20553 11655 20587
rect 14565 20553 14599 20587
rect 15577 20553 15611 20587
rect 16681 20553 16715 20587
rect 17693 20553 17727 20587
rect 19809 20553 19843 20587
rect 1501 20485 1535 20519
rect 3157 20485 3191 20519
rect 6561 20485 6595 20519
rect 14105 20485 14139 20519
rect 18613 20485 18647 20519
rect 20453 20485 20487 20519
rect 2237 20417 2271 20451
rect 2881 20417 2915 20451
rect 3893 20417 3927 20451
rect 4629 20417 4663 20451
rect 5449 20439 5483 20473
rect 5541 20417 5575 20451
rect 5718 20417 5752 20451
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 6653 20417 6687 20451
rect 6745 20417 6779 20451
rect 7665 20417 7699 20451
rect 7849 20417 7883 20451
rect 7941 20417 7975 20451
rect 8217 20417 8251 20451
rect 8677 20417 8711 20451
rect 8861 20417 8895 20451
rect 8953 20417 8987 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10149 20417 10183 20451
rect 10609 20417 10643 20451
rect 11621 20417 11655 20451
rect 11805 20417 11839 20451
rect 11897 20417 11931 20451
rect 12173 20417 12207 20451
rect 12725 20417 12759 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 13277 20417 13311 20451
rect 13921 20417 13955 20451
rect 14749 20417 14783 20451
rect 14841 20417 14875 20451
rect 15117 20417 15151 20451
rect 15761 20417 15795 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 16957 20417 16991 20451
rect 17233 20417 17267 20451
rect 17877 20417 17911 20451
rect 18797 20417 18831 20451
rect 19717 20417 19751 20451
rect 1685 20349 1719 20383
rect 3157 20349 3191 20383
rect 4169 20349 4203 20383
rect 10701 20349 10735 20383
rect 18153 20349 18187 20383
rect 6929 20281 6963 20315
rect 8033 20281 8067 20315
rect 13185 20281 13219 20315
rect 18061 20281 18095 20315
rect 2973 20213 3007 20247
rect 4077 20213 4111 20247
rect 4721 20213 4755 20247
rect 5273 20213 5307 20247
rect 8125 20213 8159 20247
rect 9137 20213 9171 20247
rect 9689 20213 9723 20247
rect 10609 20213 10643 20247
rect 12081 20213 12115 20247
rect 15025 20213 15059 20247
rect 16037 20213 16071 20247
rect 17141 20213 17175 20247
rect 18981 20213 19015 20247
rect 20545 20213 20579 20247
rect 6469 20009 6503 20043
rect 7021 20009 7055 20043
rect 10885 20009 10919 20043
rect 13369 20009 13403 20043
rect 15761 20009 15795 20043
rect 16405 20009 16439 20043
rect 17141 20009 17175 20043
rect 18613 20009 18647 20043
rect 3801 19941 3835 19975
rect 9505 19941 9539 19975
rect 14749 19941 14783 19975
rect 17969 19941 18003 19975
rect 4353 19873 4387 19907
rect 7389 19873 7423 19907
rect 7481 19873 7515 19907
rect 8309 19873 8343 19907
rect 9965 19873 9999 19907
rect 10149 19873 10183 19907
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 5457 19805 5491 19839
rect 5641 19805 5675 19839
rect 7297 19805 7331 19839
rect 7573 19805 7607 19839
rect 7757 19805 7791 19839
rect 8217 19805 8251 19839
rect 11437 19805 11471 19839
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 13277 19805 13311 19839
rect 15669 19805 15703 19839
rect 16313 19805 16347 19839
rect 17785 19805 17819 19839
rect 20453 19805 20487 19839
rect 2881 19737 2915 19771
rect 3065 19737 3099 19771
rect 6377 19737 6411 19771
rect 10793 19737 10827 19771
rect 14565 19737 14599 19771
rect 17049 19737 17083 19771
rect 18521 19737 18555 19771
rect 19809 19737 19843 19771
rect 3249 19669 3283 19703
rect 4169 19669 4203 19703
rect 4261 19669 4295 19703
rect 5825 19669 5859 19703
rect 9873 19669 9907 19703
rect 11529 19669 11563 19703
rect 12357 19669 12391 19703
rect 12725 19669 12759 19703
rect 19901 19669 19935 19703
rect 20637 19669 20671 19703
rect 1593 19465 1627 19499
rect 2973 19465 3007 19499
rect 4077 19465 4111 19499
rect 5089 19465 5123 19499
rect 9045 19465 9079 19499
rect 13093 19465 13127 19499
rect 20637 19465 20671 19499
rect 6745 19397 6779 19431
rect 8401 19397 8435 19431
rect 12173 19397 12207 19431
rect 12265 19397 12299 19431
rect 14013 19397 14047 19431
rect 19809 19397 19843 19431
rect 1501 19329 1535 19363
rect 2145 19329 2179 19363
rect 2329 19329 2363 19363
rect 3433 19329 3467 19363
rect 4261 19329 4295 19363
rect 4537 19329 4571 19363
rect 4997 19329 5031 19363
rect 5641 19329 5675 19363
rect 6653 19329 6687 19363
rect 6837 19329 6871 19363
rect 7113 19329 7147 19363
rect 7665 19329 7699 19363
rect 8309 19329 8343 19363
rect 9229 19329 9263 19363
rect 9413 19329 9447 19363
rect 9505 19329 9539 19363
rect 9965 19329 9999 19363
rect 10149 19329 10183 19363
rect 10241 19329 10275 19363
rect 10517 19329 10551 19363
rect 11989 19329 12023 19363
rect 12357 19329 12391 19363
rect 13001 19329 13035 19363
rect 14105 19329 14139 19363
rect 14841 19329 14875 19363
rect 15761 19329 15795 19363
rect 15853 19329 15887 19363
rect 16037 19329 16071 19363
rect 16129 19329 16163 19363
rect 16681 19329 16715 19363
rect 17785 19329 17819 19363
rect 17877 19329 17911 19363
rect 19073 19329 19107 19363
rect 20545 19329 20579 19363
rect 2513 19261 2547 19295
rect 3341 19261 3375 19295
rect 10425 19261 10459 19295
rect 13921 19261 13955 19295
rect 14289 19261 14323 19295
rect 14381 19261 14415 19295
rect 18061 19261 18095 19295
rect 19993 19261 20027 19295
rect 3617 19193 3651 19227
rect 6377 19193 6411 19227
rect 12541 19193 12575 19227
rect 14105 19193 14139 19227
rect 19257 19193 19291 19227
rect 4445 19125 4479 19159
rect 5733 19125 5767 19159
rect 7021 19125 7055 19159
rect 7757 19125 7791 19159
rect 10333 19125 10367 19159
rect 14933 19125 14967 19159
rect 15577 19125 15611 19159
rect 16773 19125 16807 19159
rect 17969 19125 18003 19159
rect 1593 18921 1627 18955
rect 2881 18921 2915 18955
rect 3893 18921 3927 18955
rect 5365 18921 5399 18955
rect 5825 18921 5859 18955
rect 8217 18921 8251 18955
rect 11345 18921 11379 18955
rect 14197 18921 14231 18955
rect 16773 18921 16807 18955
rect 18613 18921 18647 18955
rect 19625 18921 19659 18955
rect 9873 18853 9907 18887
rect 11897 18853 11931 18887
rect 12541 18853 12575 18887
rect 17325 18853 17359 18887
rect 2237 18785 2271 18819
rect 5549 18785 5583 18819
rect 10517 18785 10551 18819
rect 13185 18785 13219 18819
rect 17877 18785 17911 18819
rect 20269 18785 20303 18819
rect 1961 18717 1995 18751
rect 2789 18717 2823 18751
rect 3801 18717 3835 18751
rect 4721 18717 4755 18751
rect 5641 18717 5675 18751
rect 6469 18717 6503 18751
rect 6929 18717 6963 18751
rect 8401 18717 8435 18751
rect 9045 18717 9079 18751
rect 10241 18717 10275 18751
rect 11470 18717 11504 18751
rect 11989 18717 12023 18751
rect 12909 18717 12943 18751
rect 14105 18717 14139 18751
rect 14381 18717 14415 18751
rect 14565 18717 14599 18751
rect 15485 18717 15519 18751
rect 15577 18717 15611 18751
rect 15669 18717 15703 18751
rect 15853 18717 15887 18751
rect 16497 18717 16531 18751
rect 16589 18717 16623 18751
rect 16865 18717 16899 18751
rect 17785 18717 17819 18751
rect 18521 18717 18555 18751
rect 5365 18649 5399 18683
rect 16313 18649 16347 18683
rect 20085 18649 20119 18683
rect 2053 18581 2087 18615
rect 4813 18581 4847 18615
rect 6285 18581 6319 18615
rect 7113 18581 7147 18615
rect 9137 18581 9171 18615
rect 10333 18581 10367 18615
rect 11529 18581 11563 18615
rect 13001 18581 13035 18615
rect 14749 18581 14783 18615
rect 15209 18581 15243 18615
rect 17693 18581 17727 18615
rect 19993 18581 20027 18615
rect 1685 18377 1719 18411
rect 2605 18377 2639 18411
rect 3433 18377 3467 18411
rect 3525 18377 3559 18411
rect 5825 18377 5859 18411
rect 7021 18377 7055 18411
rect 11529 18377 11563 18411
rect 12541 18377 12575 18411
rect 14381 18377 14415 18411
rect 17141 18377 17175 18411
rect 19809 18377 19843 18411
rect 19993 18377 20027 18411
rect 2421 18309 2455 18343
rect 5549 18309 5583 18343
rect 6745 18309 6779 18343
rect 7941 18309 7975 18343
rect 10609 18309 10643 18343
rect 1593 18241 1627 18275
rect 2237 18241 2271 18275
rect 3249 18241 3283 18275
rect 4077 18241 4111 18275
rect 5273 18241 5307 18275
rect 5457 18241 5491 18275
rect 5641 18241 5675 18275
rect 6377 18241 6411 18275
rect 6470 18241 6504 18275
rect 6653 18241 6687 18275
rect 6842 18241 6876 18275
rect 7849 18241 7883 18275
rect 8309 18241 8343 18275
rect 8677 18241 8711 18275
rect 8861 18241 8895 18275
rect 9689 18241 9723 18275
rect 10517 18241 10551 18275
rect 11713 18241 11747 18275
rect 11805 18241 11839 18275
rect 12081 18241 12115 18275
rect 12725 18241 12759 18275
rect 12817 18241 12851 18275
rect 13093 18241 13127 18275
rect 13553 18241 13587 18275
rect 14289 18241 14323 18275
rect 15945 18241 15979 18275
rect 16129 18241 16163 18275
rect 17325 18241 17359 18275
rect 17601 18241 17635 18275
rect 18153 18241 18187 18275
rect 19073 18241 19107 18275
rect 19990 18241 20024 18275
rect 20453 18241 20487 18275
rect 3065 18173 3099 18207
rect 3617 18173 3651 18207
rect 8401 18173 8435 18207
rect 9781 18173 9815 18207
rect 9965 18173 9999 18207
rect 13645 18173 13679 18207
rect 15669 18173 15703 18207
rect 11989 18105 12023 18139
rect 4169 18037 4203 18071
rect 9321 18037 9355 18071
rect 13001 18037 13035 18071
rect 15393 18037 15427 18071
rect 15761 18037 15795 18071
rect 15853 18037 15887 18071
rect 17509 18037 17543 18071
rect 18245 18037 18279 18071
rect 19257 18037 19291 18071
rect 20361 18037 20395 18071
rect 5457 17833 5491 17867
rect 6469 17833 6503 17867
rect 7389 17833 7423 17867
rect 7941 17833 7975 17867
rect 12081 17833 12115 17867
rect 12725 17833 12759 17867
rect 13369 17833 13403 17867
rect 14473 17833 14507 17867
rect 15117 17833 15151 17867
rect 15669 17833 15703 17867
rect 16773 17833 16807 17867
rect 18521 17833 18555 17867
rect 8953 17765 8987 17799
rect 9965 17765 9999 17799
rect 11529 17765 11563 17799
rect 18613 17765 18647 17799
rect 19993 17765 20027 17799
rect 20545 17765 20579 17799
rect 4353 17697 4387 17731
rect 8401 17697 8435 17731
rect 9413 17697 9447 17731
rect 10241 17697 10275 17731
rect 14105 17697 14139 17731
rect 16129 17697 16163 17731
rect 2973 17629 3007 17663
rect 3157 17629 3191 17663
rect 3249 17629 3283 17663
rect 5273 17629 5307 17663
rect 5549 17629 5583 17663
rect 6193 17629 6227 17663
rect 6377 17629 6411 17663
rect 6561 17629 6595 17663
rect 7021 17629 7055 17663
rect 7205 17629 7239 17663
rect 8125 17629 8159 17663
rect 8309 17629 8343 17663
rect 9045 17629 9079 17663
rect 9229 17629 9263 17663
rect 9505 17629 9539 17663
rect 10057 17629 10091 17663
rect 10425 17629 10459 17663
rect 10517 17629 10551 17663
rect 11345 17629 11379 17663
rect 11989 17629 12023 17663
rect 12633 17629 12667 17663
rect 13553 17629 13587 17663
rect 14289 17629 14323 17663
rect 14565 17629 14599 17663
rect 15025 17629 15059 17663
rect 15669 17629 15703 17663
rect 15853 17629 15887 17663
rect 15945 17629 15979 17663
rect 16221 17629 16255 17663
rect 16681 17629 16715 17663
rect 17325 17629 17359 17663
rect 18153 17629 18187 17663
rect 18337 17629 18371 17663
rect 18429 17629 18463 17663
rect 18705 17629 18739 17663
rect 19566 17629 19600 17663
rect 20085 17629 20119 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 1869 17561 1903 17595
rect 2789 17561 2823 17595
rect 4261 17561 4295 17595
rect 17509 17561 17543 17595
rect 1961 17493 1995 17527
rect 3801 17493 3835 17527
rect 4169 17493 4203 17527
rect 5089 17493 5123 17527
rect 9137 17493 9171 17527
rect 10149 17493 10183 17527
rect 17693 17493 17727 17527
rect 19441 17493 19475 17527
rect 19625 17493 19659 17527
rect 1777 17289 1811 17323
rect 2513 17289 2547 17323
rect 3617 17289 3651 17323
rect 5273 17289 5307 17323
rect 6561 17289 6595 17323
rect 8953 17289 8987 17323
rect 13921 17289 13955 17323
rect 14381 17289 14415 17323
rect 20269 17289 20303 17323
rect 20637 17289 20671 17323
rect 1961 17153 1995 17187
rect 2697 17153 2731 17187
rect 3801 17153 3835 17187
rect 4077 17153 4111 17187
rect 5270 17153 5304 17187
rect 5641 17153 5675 17187
rect 6377 17153 6411 17187
rect 6561 17153 6595 17187
rect 7021 17153 7055 17187
rect 7205 17153 7239 17187
rect 7297 17153 7331 17187
rect 7573 17153 7607 17187
rect 8677 17153 8711 17187
rect 9413 17153 9447 17187
rect 10057 17153 10091 17187
rect 10701 17153 10735 17187
rect 11713 17153 11747 17187
rect 12173 17153 12207 17187
rect 12909 17153 12943 17187
rect 14289 17153 14323 17187
rect 15393 17153 15427 17187
rect 15577 17153 15611 17187
rect 15669 17153 15703 17187
rect 17325 17153 17359 17187
rect 17417 17153 17451 17187
rect 17693 17153 17727 17187
rect 18429 17153 18463 17187
rect 18613 17153 18647 17187
rect 19533 17153 19567 17187
rect 20453 17153 20487 17187
rect 20729 17153 20763 17187
rect 5733 17085 5767 17119
rect 8953 17085 8987 17119
rect 14473 17085 14507 17119
rect 17233 17085 17267 17119
rect 19809 17085 19843 17119
rect 3985 17017 4019 17051
rect 8769 17017 8803 17051
rect 17417 17017 17451 17051
rect 18797 17017 18831 17051
rect 5089 16949 5123 16983
rect 7021 16949 7055 16983
rect 7481 16949 7515 16983
rect 9597 16949 9631 16983
rect 10241 16949 10275 16983
rect 10793 16949 10827 16983
rect 11529 16949 11563 16983
rect 12357 16949 12391 16983
rect 13001 16949 13035 16983
rect 15485 16949 15519 16983
rect 15853 16949 15887 16983
rect 17601 16949 17635 16983
rect 19349 16949 19383 16983
rect 19717 16949 19751 16983
rect 3617 16745 3651 16779
rect 5273 16745 5307 16779
rect 7113 16745 7147 16779
rect 14381 16745 14415 16779
rect 15577 16745 15611 16779
rect 16037 16745 16071 16779
rect 19441 16745 19475 16779
rect 2053 16541 2087 16575
rect 2513 16541 2547 16575
rect 3985 16677 4019 16711
rect 7297 16677 7331 16711
rect 5365 16609 5399 16643
rect 10425 16609 10459 16643
rect 14105 16609 14139 16643
rect 14657 16609 14691 16643
rect 17693 16609 17727 16643
rect 18245 16609 18279 16643
rect 19901 16609 19935 16643
rect 20085 16609 20119 16643
rect 3801 16541 3835 16575
rect 4445 16541 4479 16575
rect 5089 16541 5123 16575
rect 5181 16541 5215 16575
rect 5917 16541 5951 16575
rect 6837 16541 6871 16575
rect 7205 16541 7239 16575
rect 7573 16541 7607 16575
rect 11529 16541 11563 16575
rect 12909 16541 12943 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 14519 16541 14553 16575
rect 15577 16541 15611 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 16129 16541 16163 16575
rect 16957 16541 16991 16575
rect 17417 16541 17451 16575
rect 17509 16541 17543 16575
rect 18429 16541 18463 16575
rect 18705 16541 18739 16575
rect 19809 16541 19843 16575
rect 3617 16473 3651 16507
rect 1869 16405 1903 16439
rect 2697 16405 2731 16439
rect 4629 16405 4663 16439
rect 6009 16405 6043 16439
rect 7481 16405 7515 16439
rect 9781 16405 9815 16439
rect 10149 16405 10183 16439
rect 10241 16405 10275 16439
rect 11713 16405 11747 16439
rect 12725 16405 12759 16439
rect 13369 16405 13403 16439
rect 16773 16405 16807 16439
rect 17693 16405 17727 16439
rect 18613 16405 18647 16439
rect 1593 16201 1627 16235
rect 4353 16201 4387 16235
rect 5089 16201 5123 16235
rect 7113 16201 7147 16235
rect 12173 16201 12207 16235
rect 13461 16201 13495 16235
rect 15393 16201 15427 16235
rect 17693 16201 17727 16235
rect 1961 16133 1995 16167
rect 7205 16133 7239 16167
rect 12265 16133 12299 16167
rect 19165 16133 19199 16167
rect 3341 16065 3375 16099
rect 3617 16065 3651 16099
rect 4169 16065 4203 16099
rect 4813 16065 4847 16099
rect 5549 16065 5583 16099
rect 5733 16065 5767 16099
rect 10333 16065 10367 16099
rect 10517 16065 10551 16099
rect 11989 16065 12023 16099
rect 12817 16065 12851 16099
rect 13461 16065 13495 16099
rect 14565 16065 14599 16099
rect 14657 16065 14691 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 15853 16065 15887 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 16681 16065 16715 16099
rect 20177 16065 20211 16099
rect 2053 15997 2087 16031
rect 2237 15997 2271 16031
rect 3249 15997 3283 16031
rect 3709 15997 3743 16031
rect 5089 15997 5123 16031
rect 7297 15997 7331 16031
rect 10057 15997 10091 16031
rect 11805 15997 11839 16031
rect 12357 15997 12391 16031
rect 13737 15997 13771 16031
rect 17785 15997 17819 16031
rect 17877 15997 17911 16031
rect 19809 15997 19843 16031
rect 20269 15997 20303 16031
rect 4905 15929 4939 15963
rect 5549 15929 5583 15963
rect 10149 15929 10183 15963
rect 13553 15929 13587 15963
rect 16773 15929 16807 15963
rect 19349 15929 19383 15963
rect 3065 15861 3099 15895
rect 6745 15861 6779 15895
rect 9781 15861 9815 15895
rect 10241 15861 10275 15895
rect 12909 15861 12943 15895
rect 14381 15861 14415 15895
rect 14841 15861 14875 15895
rect 15761 15861 15795 15895
rect 17325 15861 17359 15895
rect 20453 15861 20487 15895
rect 2697 15657 2731 15691
rect 5365 15657 5399 15691
rect 8953 15657 8987 15691
rect 9873 15657 9907 15691
rect 15945 15657 15979 15691
rect 17049 15657 17083 15691
rect 17601 15657 17635 15691
rect 18613 15657 18647 15691
rect 12449 15589 12483 15623
rect 13093 15589 13127 15623
rect 3157 15521 3191 15555
rect 4813 15521 4847 15555
rect 5825 15521 5859 15555
rect 5917 15521 5951 15555
rect 7481 15521 7515 15555
rect 7665 15521 7699 15555
rect 9137 15521 9171 15555
rect 10333 15521 10367 15555
rect 11345 15521 11379 15555
rect 13277 15521 13311 15555
rect 1409 15453 1443 15487
rect 1685 15453 1719 15487
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 3249 15453 3283 15487
rect 6561 15453 6595 15487
rect 6653 15453 6687 15487
rect 7389 15453 7423 15487
rect 9229 15453 9263 15487
rect 9873 15453 9907 15487
rect 10057 15453 10091 15487
rect 10149 15453 10183 15487
rect 10425 15453 10459 15487
rect 11069 15453 11103 15487
rect 11161 15453 11195 15487
rect 11437 15453 11471 15487
rect 11897 15453 11931 15487
rect 12265 15453 12299 15487
rect 13185 15453 13219 15487
rect 14381 15453 14415 15487
rect 15393 15453 15427 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16957 15453 16991 15487
rect 17877 15453 17911 15487
rect 18521 15453 18555 15487
rect 19257 15453 19291 15487
rect 19901 15453 19935 15487
rect 20177 15453 20211 15487
rect 4537 15385 4571 15419
rect 7665 15385 7699 15419
rect 8953 15385 8987 15419
rect 12081 15385 12115 15419
rect 12173 15385 12207 15419
rect 12909 15385 12943 15419
rect 15669 15385 15703 15419
rect 17601 15385 17635 15419
rect 4169 15317 4203 15351
rect 4629 15317 4663 15351
rect 5733 15317 5767 15351
rect 9413 15317 9447 15351
rect 10885 15317 10919 15351
rect 13001 15317 13035 15351
rect 14473 15317 14507 15351
rect 17785 15317 17819 15351
rect 19349 15317 19383 15351
rect 2145 15113 2179 15147
rect 4629 15113 4663 15147
rect 5365 15113 5399 15147
rect 7573 15113 7607 15147
rect 12449 15113 12483 15147
rect 20177 15113 20211 15147
rect 3249 15045 3283 15079
rect 4445 15045 4479 15079
rect 10057 15045 10091 15079
rect 10149 15045 10183 15079
rect 12541 15045 12575 15079
rect 2053 14977 2087 15011
rect 2973 14977 3007 15011
rect 4721 14977 4755 15011
rect 5549 14977 5583 15011
rect 5825 14977 5859 15011
rect 7665 14977 7699 15011
rect 10701 14977 10735 15011
rect 12081 14977 12115 15011
rect 12633 14977 12667 15011
rect 13461 14977 13495 15011
rect 14105 14977 14139 15011
rect 14381 14977 14415 15011
rect 14657 14977 14691 15011
rect 14841 14977 14875 15011
rect 15761 14977 15795 15011
rect 15853 14977 15887 15011
rect 15945 14977 15979 15011
rect 16129 14977 16163 15011
rect 16681 14977 16715 15011
rect 17877 14977 17911 15011
rect 18061 14977 18095 15011
rect 19073 14977 19107 15011
rect 20085 14977 20119 15011
rect 2881 14909 2915 14943
rect 3341 14909 3375 14943
rect 7297 14909 7331 14943
rect 9965 14909 9999 14943
rect 11897 14909 11931 14943
rect 12340 14909 12374 14943
rect 14473 14909 14507 14943
rect 16773 14909 16807 14943
rect 20269 14909 20303 14943
rect 4445 14841 4479 14875
rect 7205 14841 7239 14875
rect 9597 14841 9631 14875
rect 19257 14841 19291 14875
rect 2697 14773 2731 14807
rect 5733 14773 5767 14807
rect 6929 14773 6963 14807
rect 7389 14773 7423 14807
rect 10793 14773 10827 14807
rect 13553 14773 13587 14807
rect 15485 14773 15519 14807
rect 17877 14773 17911 14807
rect 19717 14773 19751 14807
rect 2789 14569 2823 14603
rect 4905 14569 4939 14603
rect 5273 14569 5307 14603
rect 5825 14569 5859 14603
rect 6929 14569 6963 14603
rect 9689 14569 9723 14603
rect 10609 14569 10643 14603
rect 12449 14569 12483 14603
rect 14105 14569 14139 14603
rect 14565 14569 14599 14603
rect 16405 14569 16439 14603
rect 17141 14569 17175 14603
rect 17877 14569 17911 14603
rect 19441 14569 19475 14603
rect 20729 14569 20763 14603
rect 2329 14501 2363 14535
rect 10977 14501 11011 14535
rect 12909 14501 12943 14535
rect 13185 14501 13219 14535
rect 18245 14501 18279 14535
rect 7205 14433 7239 14467
rect 7573 14433 7607 14467
rect 10701 14433 10735 14467
rect 13369 14433 13403 14467
rect 17325 14433 17359 14467
rect 19901 14433 19935 14467
rect 2513 14365 2547 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 3801 14365 3835 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 5733 14365 5767 14399
rect 6837 14365 6871 14399
rect 7297 14365 7331 14399
rect 7665 14365 7699 14399
rect 9045 14365 9079 14399
rect 9229 14365 9263 14399
rect 9873 14365 9907 14399
rect 10057 14365 10091 14399
rect 10149 14365 10183 14399
rect 10609 14365 10643 14399
rect 11805 14365 11839 14399
rect 11953 14365 11987 14399
rect 12289 14365 12323 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 13553 14365 13587 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 14657 14365 14691 14399
rect 15117 14365 15151 14399
rect 16589 14365 16623 14399
rect 17049 14365 17083 14399
rect 17877 14365 17911 14399
rect 17969 14365 18003 14399
rect 19625 14365 19659 14399
rect 19809 14365 19843 14399
rect 20545 14365 20579 14399
rect 1685 14297 1719 14331
rect 1869 14297 1903 14331
rect 9137 14297 9171 14331
rect 12081 14297 12115 14331
rect 12173 14297 12207 14331
rect 20361 14297 20395 14331
rect 3893 14229 3927 14263
rect 15209 14229 15243 14263
rect 17325 14229 17359 14263
rect 21557 14229 21591 14263
rect 3341 14025 3375 14059
rect 5549 14025 5583 14059
rect 6837 14025 6871 14059
rect 7481 14025 7515 14059
rect 9689 14025 9723 14059
rect 11897 14025 11931 14059
rect 14111 14025 14145 14059
rect 16681 14025 16715 14059
rect 17141 14025 17175 14059
rect 18061 14025 18095 14059
rect 19993 14025 20027 14059
rect 20177 14025 20211 14059
rect 4537 13957 4571 13991
rect 6745 13957 6779 13991
rect 8125 13957 8159 13991
rect 12817 13957 12851 13991
rect 14197 13957 14231 13991
rect 1501 13889 1535 13923
rect 2329 13889 2363 13923
rect 2421 13889 2455 13923
rect 2697 13889 2731 13923
rect 3157 13889 3191 13923
rect 3433 13889 3467 13923
rect 4445 13889 4479 13923
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 2605 13821 2639 13855
rect 5273 13821 5307 13855
rect 7573 13889 7607 13923
rect 8033 13889 8067 13923
rect 9873 13889 9907 13923
rect 10149 13889 10183 13923
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 11894 13889 11928 13923
rect 12357 13889 12391 13923
rect 13001 13889 13035 13923
rect 14013 13889 14047 13923
rect 14289 13889 14323 13923
rect 14749 13889 14783 13923
rect 14933 13889 14967 13923
rect 17049 13889 17083 13923
rect 17877 13889 17911 13923
rect 18889 13889 18923 13923
rect 19073 13889 19107 13923
rect 19165 13889 19199 13923
rect 19441 13889 19475 13923
rect 20174 13889 20208 13923
rect 20545 13889 20579 13923
rect 10885 13821 10919 13855
rect 12265 13821 12299 13855
rect 13185 13821 13219 13855
rect 17325 13821 17359 13855
rect 17969 13821 18003 13855
rect 18153 13821 18187 13855
rect 18429 13821 18463 13855
rect 20637 13821 20671 13855
rect 6745 13753 6779 13787
rect 7205 13753 7239 13787
rect 7297 13753 7331 13787
rect 10057 13753 10091 13787
rect 14749 13753 14783 13787
rect 19257 13753 19291 13787
rect 1593 13685 1627 13719
rect 2145 13685 2179 13719
rect 3157 13685 3191 13719
rect 5181 13685 5215 13719
rect 7113 13685 7147 13719
rect 10793 13685 10827 13719
rect 11713 13685 11747 13719
rect 18337 13685 18371 13719
rect 19349 13685 19383 13719
rect 2881 13481 2915 13515
rect 3893 13481 3927 13515
rect 5733 13481 5767 13515
rect 12449 13481 12483 13515
rect 14197 13481 14231 13515
rect 14933 13481 14967 13515
rect 15945 13481 15979 13515
rect 16957 13481 16991 13515
rect 17785 13481 17819 13515
rect 15209 13413 15243 13447
rect 17141 13413 17175 13447
rect 19257 13413 19291 13447
rect 2145 13345 2179 13379
rect 2237 13345 2271 13379
rect 7113 13345 7147 13379
rect 9045 13345 9079 13379
rect 9229 13345 9263 13379
rect 9321 13345 9355 13379
rect 10517 13345 10551 13379
rect 11805 13345 11839 13379
rect 14841 13345 14875 13379
rect 15761 13345 15795 13379
rect 16589 13345 16623 13379
rect 16773 13345 16807 13379
rect 18705 13345 18739 13379
rect 19901 13345 19935 13379
rect 2881 13277 2915 13311
rect 3065 13277 3099 13311
rect 3801 13277 3835 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 6653 13277 6687 13311
rect 6837 13277 6871 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 9505 13277 9539 13311
rect 10425 13277 10459 13311
rect 11161 13277 11195 13311
rect 12173 13277 12207 13311
rect 12265 13277 12299 13311
rect 14105 13277 14139 13311
rect 14749 13277 14783 13311
rect 15025 13277 15059 13311
rect 15945 13277 15979 13311
rect 2053 13209 2087 13243
rect 5365 13209 5399 13243
rect 5549 13209 5583 13243
rect 15669 13209 15703 13243
rect 16957 13277 16991 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 19625 13277 19659 13311
rect 16681 13209 16715 13243
rect 18521 13209 18555 13243
rect 20545 13209 20579 13243
rect 1685 13141 1719 13175
rect 4813 13141 4847 13175
rect 6653 13141 6687 13175
rect 9045 13141 9079 13175
rect 9137 13141 9171 13175
rect 9965 13141 9999 13175
rect 10333 13141 10367 13175
rect 11253 13141 11287 13175
rect 16129 13141 16163 13175
rect 16589 13141 16623 13175
rect 19717 13141 19751 13175
rect 20637 13141 20671 13175
rect 1961 12937 1995 12971
rect 10241 12937 10275 12971
rect 11989 12937 12023 12971
rect 13277 12937 13311 12971
rect 14657 12937 14691 12971
rect 16681 12937 16715 12971
rect 19441 12937 19475 12971
rect 19625 12937 19659 12971
rect 3801 12869 3835 12903
rect 5273 12869 5307 12903
rect 7481 12869 7515 12903
rect 1869 12801 1903 12835
rect 2881 12801 2915 12835
rect 2973 12801 3007 12835
rect 3249 12801 3283 12835
rect 3709 12801 3743 12835
rect 5089 12801 5123 12835
rect 5365 12801 5399 12835
rect 6837 12801 6871 12835
rect 7665 12801 7699 12835
rect 7757 12801 7791 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10425 12801 10459 12835
rect 11897 12801 11931 12835
rect 13185 12801 13219 12835
rect 14289 12801 14323 12835
rect 14749 12801 14783 12835
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 17601 12801 17635 12835
rect 18613 12801 18647 12835
rect 19622 12801 19656 12835
rect 20085 12801 20119 12835
rect 20545 12801 20579 12835
rect 3157 12733 3191 12767
rect 9321 12733 9355 12767
rect 10701 12733 10735 12767
rect 12173 12733 12207 12767
rect 13369 12733 13403 12767
rect 14473 12733 14507 12767
rect 17141 12733 17175 12767
rect 17693 12733 17727 12767
rect 9689 12665 9723 12699
rect 16129 12665 16163 12699
rect 2697 12597 2731 12631
rect 4905 12597 4939 12631
rect 6929 12597 6963 12631
rect 7481 12597 7515 12631
rect 7941 12597 7975 12631
rect 10609 12597 10643 12631
rect 11529 12597 11563 12631
rect 12817 12597 12851 12631
rect 14013 12597 14047 12631
rect 14381 12597 14415 12631
rect 17049 12597 17083 12631
rect 18705 12597 18739 12631
rect 19993 12597 20027 12631
rect 20637 12597 20671 12631
rect 1409 12393 1443 12427
rect 3157 12393 3191 12427
rect 6837 12393 6871 12427
rect 11713 12393 11747 12427
rect 12449 12393 12483 12427
rect 13461 12393 13495 12427
rect 14105 12393 14139 12427
rect 15301 12393 15335 12427
rect 17601 12393 17635 12427
rect 20085 12393 20119 12427
rect 2881 12325 2915 12359
rect 6193 12325 6227 12359
rect 10241 12325 10275 12359
rect 2973 12257 3007 12291
rect 3249 12257 3283 12291
rect 5089 12257 5123 12291
rect 5273 12257 5307 12291
rect 7021 12257 7055 12291
rect 7941 12257 7975 12291
rect 14565 12257 14599 12291
rect 1593 12189 1627 12223
rect 2053 12189 2087 12223
rect 2789 12189 2823 12223
rect 6009 12189 6043 12223
rect 6285 12189 6319 12223
rect 6745 12189 6779 12223
rect 7481 12189 7515 12223
rect 7665 12189 7699 12223
rect 7757 12189 7791 12223
rect 8033 12189 8067 12223
rect 10057 12189 10091 12223
rect 10818 12189 10852 12223
rect 11529 12189 11563 12223
rect 12265 12189 12299 12223
rect 13369 12189 13403 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 14381 12189 14415 12223
rect 14657 12189 14691 12223
rect 15117 12189 15151 12223
rect 15853 12189 15887 12223
rect 16681 12189 16715 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 17693 12189 17727 12223
rect 18153 12189 18187 12223
rect 20269 12189 20303 12223
rect 20545 12189 20579 12223
rect 4997 12121 5031 12155
rect 5825 12121 5859 12155
rect 19441 12121 19475 12155
rect 20453 12121 20487 12155
rect 2145 12053 2179 12087
rect 2881 12053 2915 12087
rect 4629 12053 4663 12087
rect 7021 12053 7055 12087
rect 7481 12053 7515 12087
rect 10977 12053 11011 12087
rect 16037 12053 16071 12087
rect 16497 12053 16531 12087
rect 17141 12053 17175 12087
rect 18245 12053 18279 12087
rect 19533 12053 19567 12087
rect 2329 11849 2363 11883
rect 4905 11849 4939 11883
rect 5365 11849 5399 11883
rect 8309 11849 8343 11883
rect 11713 11849 11747 11883
rect 14841 11849 14875 11883
rect 15393 11849 15427 11883
rect 16865 11849 16899 11883
rect 19073 11849 19107 11883
rect 9229 11781 9263 11815
rect 9873 11781 9907 11815
rect 20269 11781 20303 11815
rect 20453 11781 20487 11815
rect 1501 11713 1535 11747
rect 2326 11713 2360 11747
rect 2697 11713 2731 11747
rect 2789 11713 2823 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 4261 11713 4295 11747
rect 5273 11713 5307 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 10563 11713 10597 11747
rect 10701 11713 10735 11747
rect 11529 11713 11563 11747
rect 12265 11713 12299 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 13277 11713 13311 11747
rect 13553 11713 13587 11747
rect 14013 11713 14047 11747
rect 14657 11713 14691 11747
rect 15761 11713 15795 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 18245 11713 18279 11747
rect 18337 11713 18371 11747
rect 18613 11713 18647 11747
rect 19257 11713 19291 11747
rect 19349 11713 19383 11747
rect 19625 11713 19659 11747
rect 5457 11645 5491 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 8401 11645 8435 11679
rect 8585 11645 8619 11679
rect 10425 11645 10459 11679
rect 15853 11645 15887 11679
rect 16037 11645 16071 11679
rect 17141 11645 17175 11679
rect 20637 11645 20671 11679
rect 2145 11577 2179 11611
rect 17325 11577 17359 11611
rect 18521 11577 18555 11611
rect 1593 11509 1627 11543
rect 3249 11509 3283 11543
rect 3709 11509 3743 11543
rect 4353 11509 4387 11543
rect 7941 11509 7975 11543
rect 9321 11509 9355 11543
rect 12449 11509 12483 11543
rect 13001 11509 13035 11543
rect 13461 11509 13495 11543
rect 14105 11509 14139 11543
rect 17233 11509 17267 11543
rect 18061 11509 18095 11543
rect 19533 11509 19567 11543
rect 2513 11305 2547 11339
rect 3801 11305 3835 11339
rect 4261 11305 4295 11339
rect 6009 11305 6043 11339
rect 7205 11305 7239 11339
rect 9505 11305 9539 11339
rect 10333 11305 10367 11339
rect 11253 11305 11287 11339
rect 12725 11305 12759 11339
rect 13093 11305 13127 11339
rect 14841 11305 14875 11339
rect 15393 11305 15427 11339
rect 16589 11305 16623 11339
rect 6745 11237 6779 11271
rect 7665 11237 7699 11271
rect 4905 11169 4939 11203
rect 7481 11169 7515 11203
rect 7573 11169 7607 11203
rect 13185 11169 13219 11203
rect 14933 11169 14967 11203
rect 15577 11169 15611 11203
rect 15669 11169 15703 11203
rect 17601 11169 17635 11203
rect 17693 11169 17727 11203
rect 20177 11169 20211 11203
rect 1409 11101 1443 11135
rect 1501 11101 1535 11135
rect 2329 11101 2363 11135
rect 2513 11101 2547 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4353 11101 4387 11135
rect 4813 11101 4847 11135
rect 5917 11101 5951 11135
rect 6561 11101 6595 11135
rect 7941 11101 7975 11135
rect 9321 11101 9355 11135
rect 10149 11101 10183 11135
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 14657 11101 14691 11135
rect 14749 11101 14783 11135
rect 16044 11101 16078 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17509 11101 17543 11135
rect 18521 11101 18555 11135
rect 2053 11033 2087 11067
rect 18705 11033 18739 11067
rect 2697 10965 2731 10999
rect 7849 10965 7883 10999
rect 11621 10965 11655 10999
rect 15761 10965 15795 10999
rect 15945 10965 15979 10999
rect 17141 10965 17175 10999
rect 19625 10965 19659 10999
rect 19993 10965 20027 10999
rect 20085 10965 20119 10999
rect 2697 10761 2731 10795
rect 9505 10761 9539 10795
rect 14749 10761 14783 10795
rect 15853 10761 15887 10795
rect 18521 10761 18555 10795
rect 19625 10761 19659 10795
rect 2329 10693 2363 10727
rect 2421 10693 2455 10727
rect 4261 10693 4295 10727
rect 6377 10693 6411 10727
rect 12817 10693 12851 10727
rect 15485 10693 15519 10727
rect 17969 10693 18003 10727
rect 1501 10625 1535 10659
rect 2145 10625 2179 10659
rect 2513 10625 2547 10659
rect 3433 10625 3467 10659
rect 3538 10625 3572 10659
rect 3638 10625 3672 10659
rect 3801 10625 3835 10659
rect 4445 10625 4479 10659
rect 4537 10625 4571 10659
rect 4721 10625 4755 10659
rect 4813 10625 4847 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 6653 10625 6687 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7573 10625 7607 10659
rect 7757 10625 7791 10659
rect 7849 10625 7883 10659
rect 8125 10625 8159 10659
rect 8585 10625 8619 10659
rect 9321 10625 9355 10659
rect 10057 10625 10091 10659
rect 10793 10625 10827 10659
rect 11989 10625 12023 10659
rect 13829 10625 13863 10659
rect 14473 10625 14507 10659
rect 15669 10625 15703 10659
rect 16681 10625 16715 10659
rect 17877 10625 17911 10659
rect 18705 10625 18739 10659
rect 18797 10625 18831 10659
rect 19073 10625 19107 10659
rect 19809 10625 19843 10659
rect 20545 10625 20579 10659
rect 14749 10557 14783 10591
rect 18981 10557 19015 10591
rect 20085 10557 20119 10591
rect 10241 10489 10275 10523
rect 14013 10489 14047 10523
rect 1593 10421 1627 10455
rect 3157 10421 3191 10455
rect 6745 10421 6779 10455
rect 6837 10421 6871 10455
rect 7573 10421 7607 10455
rect 8033 10421 8067 10455
rect 8769 10421 8803 10455
rect 10885 10421 10919 10455
rect 14565 10421 14599 10455
rect 16773 10421 16807 10455
rect 19993 10421 20027 10455
rect 20637 10421 20671 10455
rect 2789 10217 2823 10251
rect 3985 10217 4019 10251
rect 8309 10217 8343 10251
rect 8953 10217 8987 10251
rect 10609 10217 10643 10251
rect 10701 10217 10735 10251
rect 12449 10217 12483 10251
rect 13185 10217 13219 10251
rect 16129 10217 16163 10251
rect 19349 10217 19383 10251
rect 20085 10217 20119 10251
rect 4721 10149 4755 10183
rect 10793 10149 10827 10183
rect 15485 10149 15519 10183
rect 19993 10149 20027 10183
rect 7021 10081 7055 10115
rect 9413 10081 9447 10115
rect 9597 10081 9631 10115
rect 18245 10081 18279 10115
rect 20177 10081 20211 10115
rect 2513 10013 2547 10047
rect 2605 10013 2639 10047
rect 2881 10013 2915 10047
rect 3893 10013 3927 10047
rect 4537 10013 4571 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 6837 10013 6871 10047
rect 8217 10013 8251 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11529 10013 11563 10047
rect 12265 10013 12299 10047
rect 13001 10013 13035 10047
rect 13185 10013 13219 10047
rect 15301 10013 15335 10047
rect 16037 10013 16071 10047
rect 17325 10013 17359 10047
rect 17969 10013 18003 10047
rect 18061 10013 18095 10047
rect 19257 10013 19291 10047
rect 19901 10013 19935 10047
rect 1685 9945 1719 9979
rect 2329 9945 2363 9979
rect 6929 9945 6963 9979
rect 14657 9945 14691 9979
rect 14841 9945 14875 9979
rect 17141 9945 17175 9979
rect 17509 9945 17543 9979
rect 1777 9877 1811 9911
rect 5457 9877 5491 9911
rect 6469 9877 6503 9911
rect 9321 9877 9355 9911
rect 10333 9877 10367 9911
rect 11713 9877 11747 9911
rect 13369 9877 13403 9911
rect 18245 9877 18279 9911
rect 9781 9673 9815 9707
rect 12449 9673 12483 9707
rect 13921 9673 13955 9707
rect 4721 9605 4755 9639
rect 4905 9605 4939 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 3893 9537 3927 9571
rect 4997 9537 5031 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 6377 9537 6411 9571
rect 7481 9537 7515 9571
rect 7573 9537 7607 9571
rect 11529 9537 11563 9571
rect 14473 9605 14507 9639
rect 17141 9605 17175 9639
rect 18337 9605 18371 9639
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 15117 9537 15151 9571
rect 15853 9537 15887 9571
rect 17325 9537 17359 9571
rect 18153 9537 18187 9571
rect 18429 9537 18463 9571
rect 18889 9537 18923 9571
rect 19901 9537 19935 9571
rect 20545 9537 20579 9571
rect 2605 9469 2639 9503
rect 3157 9469 3191 9503
rect 7757 9469 7791 9503
rect 8769 9469 8803 9503
rect 12449 9469 12483 9503
rect 12633 9469 12667 9503
rect 13645 9469 13679 9503
rect 18981 9469 19015 9503
rect 1501 9401 1535 9435
rect 7665 9401 7699 9435
rect 11713 9401 11747 9435
rect 17969 9401 18003 9435
rect 20361 9401 20395 9435
rect 2145 9333 2179 9367
rect 3709 9333 3743 9367
rect 4721 9333 4755 9367
rect 5549 9333 5583 9367
rect 5825 9333 5859 9367
rect 6469 9333 6503 9367
rect 12541 9333 12575 9367
rect 12909 9333 12943 9367
rect 13553 9333 13587 9367
rect 15301 9333 15335 9367
rect 16037 9333 16071 9367
rect 17509 9333 17543 9367
rect 19717 9333 19751 9367
rect 9965 9129 9999 9163
rect 15577 9129 15611 9163
rect 7389 9061 7423 9095
rect 12357 9061 12391 9095
rect 15669 9061 15703 9095
rect 4997 8993 5031 9027
rect 5181 8993 5215 9027
rect 6193 8993 6227 9027
rect 7481 8993 7515 9027
rect 15485 8993 15519 9027
rect 18153 8993 18187 9027
rect 19901 8993 19935 9027
rect 1869 8925 1903 8959
rect 2697 8925 2731 8959
rect 3801 8925 3835 8959
rect 5917 8925 5951 8959
rect 6101 8925 6135 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 8953 8925 8987 8959
rect 10149 8925 10183 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 11345 8925 11379 8959
rect 11621 8925 11655 8959
rect 12173 8925 12207 8959
rect 13001 8925 13035 8959
rect 14105 8925 14139 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 16865 8925 16899 8959
rect 17049 8925 17083 8959
rect 17141 8925 17175 8959
rect 18061 8925 18095 8959
rect 20545 8925 20579 8959
rect 4905 8857 4939 8891
rect 9045 8857 9079 8891
rect 16681 8857 16715 8891
rect 19625 8857 19659 8891
rect 20729 8857 20763 8891
rect 1961 8789 1995 8823
rect 2789 8789 2823 8823
rect 3893 8789 3927 8823
rect 4537 8789 4571 8823
rect 5733 8789 5767 8823
rect 8217 8789 8251 8823
rect 13185 8789 13219 8823
rect 14289 8789 14323 8823
rect 15209 8789 15243 8823
rect 17601 8789 17635 8823
rect 17969 8789 18003 8823
rect 19257 8789 19291 8823
rect 19717 8789 19751 8823
rect 2145 8585 2179 8619
rect 3249 8585 3283 8619
rect 4997 8585 5031 8619
rect 5365 8585 5399 8619
rect 6745 8585 6779 8619
rect 8677 8585 8711 8619
rect 8769 8585 8803 8619
rect 9321 8585 9355 8619
rect 10977 8585 11011 8619
rect 12081 8585 12115 8619
rect 14197 8585 14231 8619
rect 16957 8585 16991 8619
rect 20269 8585 20303 8619
rect 2881 8517 2915 8551
rect 5457 8517 5491 8551
rect 9965 8517 9999 8551
rect 19441 8517 19475 8551
rect 1869 8449 1903 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3065 8449 3099 8483
rect 3985 8449 4019 8483
rect 4077 8449 4111 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8493 8449 8527 8483
rect 9597 8449 9631 8483
rect 9873 8449 9907 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 12449 8449 12483 8483
rect 13277 8449 13311 8483
rect 14013 8449 14047 8483
rect 15485 8449 15519 8483
rect 17141 8449 17175 8483
rect 17877 8449 17911 8483
rect 18705 8449 18739 8483
rect 19165 8449 19199 8483
rect 19349 8449 19383 8483
rect 19533 8449 19567 8483
rect 20177 8449 20211 8483
rect 1685 8381 1719 8415
rect 2237 8381 2271 8415
rect 5549 8381 5583 8415
rect 8309 8381 8343 8415
rect 8861 8381 8895 8415
rect 9505 8381 9539 8415
rect 10701 8381 10735 8415
rect 12541 8381 12575 8415
rect 12725 8381 12759 8415
rect 15577 8381 15611 8415
rect 15761 8381 15795 8415
rect 17417 8381 17451 8415
rect 3709 8313 3743 8347
rect 7021 8313 7055 8347
rect 7113 8313 7147 8347
rect 7205 8313 7239 8347
rect 15117 8313 15151 8347
rect 17969 8313 18003 8347
rect 18521 8313 18555 8347
rect 19717 8313 19751 8347
rect 1961 8245 1995 8279
rect 10517 8245 10551 8279
rect 13461 8245 13495 8279
rect 17325 8245 17359 8279
rect 3893 8041 3927 8075
rect 5549 8041 5583 8075
rect 12909 8041 12943 8075
rect 13369 8041 13403 8075
rect 15301 8041 15335 8075
rect 16957 8041 16991 8075
rect 1869 7973 1903 8007
rect 5457 7973 5491 8007
rect 9781 7973 9815 8007
rect 11897 7973 11931 8007
rect 14749 7973 14783 8007
rect 2789 7905 2823 7939
rect 5641 7905 5675 7939
rect 7849 7905 7883 7939
rect 11989 7905 12023 7939
rect 15761 7905 15795 7939
rect 19901 7905 19935 7939
rect 1685 7837 1719 7871
rect 2513 7837 2547 7871
rect 2605 7837 2639 7871
rect 2881 7837 2915 7871
rect 3801 7837 3835 7871
rect 4445 7837 4479 7871
rect 4629 7837 4663 7871
rect 5365 7837 5399 7871
rect 6101 7837 6135 7871
rect 7665 7837 7699 7871
rect 9137 7837 9171 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 10057 7837 10091 7871
rect 10425 7837 10459 7871
rect 10609 7837 10643 7871
rect 11253 7837 11287 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13461 7837 13495 7871
rect 14565 7837 14599 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 16865 7837 16899 7871
rect 17509 7837 17543 7871
rect 17601 7837 17635 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18613 7837 18647 7871
rect 18705 7837 18739 7871
rect 19438 7837 19472 7871
rect 19809 7837 19843 7871
rect 7757 7769 7791 7803
rect 20545 7769 20579 7803
rect 2329 7701 2363 7735
rect 4537 7701 4571 7735
rect 6285 7701 6319 7735
rect 7297 7701 7331 7735
rect 8953 7701 8987 7735
rect 11069 7701 11103 7735
rect 18153 7701 18187 7735
rect 19257 7701 19291 7735
rect 19441 7701 19475 7735
rect 20637 7701 20671 7735
rect 7021 7497 7055 7531
rect 8493 7497 8527 7531
rect 9689 7497 9723 7531
rect 9873 7497 9907 7531
rect 11989 7497 12023 7531
rect 13645 7497 13679 7531
rect 18613 7497 18647 7531
rect 13461 7429 13495 7463
rect 15393 7429 15427 7463
rect 18245 7429 18279 7463
rect 19073 7429 19107 7463
rect 1869 7361 1903 7395
rect 2973 7361 3007 7395
rect 3709 7361 3743 7395
rect 3893 7361 3927 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 5457 7361 5491 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 8953 7361 8987 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 10977 7361 11011 7395
rect 11529 7361 11563 7395
rect 11805 7361 11839 7395
rect 12725 7361 12759 7395
rect 13553 7361 13587 7395
rect 14013 7361 14047 7395
rect 14933 7361 14967 7395
rect 15991 7361 16025 7395
rect 16129 7361 16163 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 17015 7361 17049 7395
rect 17233 7361 17267 7395
rect 18061 7361 18095 7395
rect 18337 7361 18371 7395
rect 18429 7361 18463 7395
rect 19257 7361 19291 7395
rect 20361 7361 20395 7395
rect 3985 7293 4019 7327
rect 8125 7293 8159 7327
rect 9781 7293 9815 7327
rect 11621 7293 11655 7327
rect 13737 7293 13771 7327
rect 15761 7293 15795 7327
rect 20453 7293 20487 7327
rect 20545 7293 20579 7327
rect 2053 7225 2087 7259
rect 5549 7225 5583 7259
rect 6653 7225 6687 7259
rect 15853 7225 15887 7259
rect 17049 7225 17083 7259
rect 3065 7157 3099 7191
rect 6377 7157 6411 7191
rect 6745 7157 6779 7191
rect 8033 7157 8067 7191
rect 9137 7157 9171 7191
rect 10149 7157 10183 7191
rect 10793 7157 10827 7191
rect 11805 7157 11839 7191
rect 12909 7157 12943 7191
rect 13921 7157 13955 7191
rect 14749 7157 14783 7191
rect 15669 7157 15703 7191
rect 17141 7157 17175 7191
rect 19441 7157 19475 7191
rect 19993 7157 20027 7191
rect 2881 6953 2915 6987
rect 16037 6953 16071 6987
rect 18613 6953 18647 6987
rect 20177 6953 20211 6987
rect 6009 6885 6043 6919
rect 7849 6885 7883 6919
rect 17601 6885 17635 6919
rect 2237 6817 2271 6851
rect 6469 6817 6503 6851
rect 7941 6817 7975 6851
rect 8217 6817 8251 6851
rect 8401 6817 8435 6851
rect 11069 6817 11103 6851
rect 12817 6817 12851 6851
rect 14933 6817 14967 6851
rect 15393 6817 15427 6851
rect 16037 6817 16071 6851
rect 18153 6817 18187 6851
rect 19901 6817 19935 6851
rect 20453 6817 20487 6851
rect 2789 6749 2823 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 4537 6749 4571 6783
rect 5365 6749 5399 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 6561 6749 6595 6783
rect 7205 6749 7239 6783
rect 8125 6749 8159 6783
rect 8953 6749 8987 6783
rect 9781 6749 9815 6783
rect 10793 6749 10827 6783
rect 10977 6749 11011 6783
rect 11897 6749 11931 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 13277 6749 13311 6783
rect 14197 6749 14231 6783
rect 15117 6749 15151 6783
rect 15301 6749 15335 6783
rect 16129 6749 16163 6783
rect 16773 6749 16807 6783
rect 17509 6749 17543 6783
rect 18337 6749 18371 6783
rect 18429 6749 18463 6783
rect 18705 6749 18739 6783
rect 19257 6749 19291 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 1961 6681 1995 6715
rect 9597 6681 9631 6715
rect 13369 6681 13403 6715
rect 15853 6681 15887 6715
rect 20361 6681 20395 6715
rect 1593 6613 1627 6647
rect 2053 6613 2087 6647
rect 3899 6613 3933 6647
rect 3985 6613 4019 6647
rect 4629 6613 4663 6647
rect 5181 6613 5215 6647
rect 7021 6613 7055 6647
rect 8033 6613 8067 6647
rect 9137 6613 9171 6647
rect 9965 6613 9999 6647
rect 10609 6613 10643 6647
rect 11989 6613 12023 6647
rect 12817 6613 12851 6647
rect 14289 6613 14323 6647
rect 14933 6613 14967 6647
rect 15025 6613 15059 6647
rect 16313 6613 16347 6647
rect 16865 6613 16899 6647
rect 19441 6613 19475 6647
rect 2053 6409 2087 6443
rect 9505 6409 9539 6443
rect 9965 6409 9999 6443
rect 10885 6409 10919 6443
rect 3341 6341 3375 6375
rect 9873 6341 9907 6375
rect 12633 6341 12667 6375
rect 14565 6341 14599 6375
rect 17785 6341 17819 6375
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2605 6273 2639 6307
rect 3065 6273 3099 6307
rect 3157 6273 3191 6307
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 4445 6273 4479 6307
rect 5089 6273 5123 6307
rect 6653 6273 6687 6307
rect 7397 6273 7431 6307
rect 8401 6273 8435 6307
rect 9045 6273 9079 6307
rect 10793 6273 10827 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 12449 6273 12483 6307
rect 13461 6273 13495 6307
rect 13645 6273 13679 6307
rect 13737 6273 13771 6307
rect 14197 6273 14231 6307
rect 14381 6273 14415 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16141 6273 16175 6307
rect 16681 6273 16715 6307
rect 18061 6273 18095 6307
rect 18153 6273 18187 6307
rect 18521 6273 18555 6307
rect 18981 6273 19015 6307
rect 19533 6273 19567 6307
rect 20545 6273 20579 6307
rect 2513 6205 2547 6239
rect 4169 6205 4203 6239
rect 4261 6205 4295 6239
rect 5365 6205 5399 6239
rect 6929 6205 6963 6239
rect 10149 6205 10183 6239
rect 16773 6205 16807 6239
rect 3065 6137 3099 6171
rect 8217 6137 8251 6171
rect 12817 6137 12851 6171
rect 15945 6137 15979 6171
rect 1409 6069 1443 6103
rect 3801 6069 3835 6103
rect 4905 6069 4939 6103
rect 5273 6069 5307 6103
rect 6469 6069 6503 6103
rect 6837 6069 6871 6103
rect 7481 6069 7515 6103
rect 8861 6069 8895 6103
rect 11529 6069 11563 6103
rect 11897 6069 11931 6103
rect 13277 6069 13311 6103
rect 16037 6069 16071 6103
rect 20637 6069 20671 6103
rect 1961 5865 1995 5899
rect 2973 5865 3007 5899
rect 4997 5865 5031 5899
rect 5917 5865 5951 5899
rect 7389 5865 7423 5899
rect 18429 5865 18463 5899
rect 18705 5865 18739 5899
rect 19441 5865 19475 5899
rect 19993 5865 20027 5899
rect 2881 5729 2915 5763
rect 3065 5729 3099 5763
rect 6469 5729 6503 5763
rect 8033 5729 8067 5763
rect 10793 5729 10827 5763
rect 12725 5729 12759 5763
rect 12909 5729 12943 5763
rect 14565 5729 14599 5763
rect 16497 5729 16531 5763
rect 18429 5729 18463 5763
rect 20545 5729 20579 5763
rect 1869 5661 1903 5695
rect 4353 5661 4387 5695
rect 4501 5661 4535 5695
rect 4818 5661 4852 5695
rect 6285 5661 6319 5695
rect 9413 5661 9447 5695
rect 9597 5661 9631 5695
rect 9689 5661 9723 5695
rect 10517 5661 10551 5695
rect 11529 5661 11563 5695
rect 11805 5661 11839 5695
rect 14289 5661 14323 5695
rect 14473 5661 14507 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 16313 5661 16347 5695
rect 16589 5661 16623 5695
rect 17601 5661 17635 5695
rect 18245 5661 18279 5695
rect 18521 5661 18555 5695
rect 19349 5661 19383 5695
rect 20453 5661 20487 5695
rect 2697 5593 2731 5627
rect 4629 5593 4663 5627
rect 4721 5593 4755 5627
rect 7849 5593 7883 5627
rect 2789 5525 2823 5559
rect 6377 5525 6411 5559
rect 7757 5525 7791 5559
rect 9229 5525 9263 5559
rect 10149 5525 10183 5559
rect 10609 5525 10643 5559
rect 11345 5525 11379 5559
rect 11713 5525 11747 5559
rect 12265 5525 12299 5559
rect 12633 5525 12667 5559
rect 14105 5525 14139 5559
rect 16129 5525 16163 5559
rect 17693 5525 17727 5559
rect 20361 5525 20395 5559
rect 5089 5321 5123 5355
rect 6653 5321 6687 5355
rect 8953 5321 8987 5355
rect 9965 5321 9999 5355
rect 10793 5321 10827 5355
rect 12173 5321 12207 5355
rect 13645 5321 13679 5355
rect 13737 5321 13771 5355
rect 16681 5321 16715 5355
rect 17049 5321 17083 5355
rect 20361 5321 20395 5355
rect 1869 5253 1903 5287
rect 9873 5253 9907 5287
rect 15945 5253 15979 5287
rect 19257 5253 19291 5287
rect 19901 5253 19935 5287
rect 20453 5253 20487 5287
rect 2053 5185 2087 5219
rect 3065 5185 3099 5219
rect 3249 5185 3283 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 5273 5185 5307 5219
rect 5365 5185 5399 5219
rect 6377 5185 6411 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 7849 5185 7883 5219
rect 8861 5185 8895 5219
rect 10701 5185 10735 5219
rect 11713 5185 11747 5219
rect 12357 5185 12391 5219
rect 12633 5185 12667 5219
rect 14473 5185 14507 5219
rect 14657 5185 14691 5219
rect 14749 5185 14783 5219
rect 15025 5185 15059 5219
rect 18061 5185 18095 5219
rect 18889 5185 18923 5219
rect 6653 5117 6687 5151
rect 10149 5117 10183 5151
rect 13829 5117 13863 5151
rect 17141 5117 17175 5151
rect 17325 5117 17359 5151
rect 18705 5117 18739 5151
rect 19993 5185 20027 5219
rect 20109 5185 20143 5219
rect 20545 5117 20579 5151
rect 4261 5049 4295 5083
rect 7665 5049 7699 5083
rect 11529 5049 11563 5083
rect 12541 5049 12575 5083
rect 16129 5049 16163 5083
rect 18889 5049 18923 5083
rect 19901 5049 19935 5083
rect 6469 4981 6503 5015
rect 7757 4981 7791 5015
rect 9505 4981 9539 5015
rect 13277 4981 13311 5015
rect 14473 4981 14507 5015
rect 14933 4981 14967 5015
rect 18153 4981 18187 5015
rect 3801 4777 3835 4811
rect 6193 4777 6227 4811
rect 9229 4777 9263 4811
rect 11345 4777 11379 4811
rect 15945 4777 15979 4811
rect 17049 4777 17083 4811
rect 18613 4777 18647 4811
rect 19901 4777 19935 4811
rect 16957 4709 16991 4743
rect 17601 4709 17635 4743
rect 1685 4641 1719 4675
rect 4445 4641 4479 4675
rect 8953 4641 8987 4675
rect 9505 4641 9539 4675
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 11805 4641 11839 4675
rect 12173 4641 12207 4675
rect 17141 4641 17175 4675
rect 1409 4573 1443 4607
rect 2881 4573 2915 4607
rect 3926 4573 3960 4607
rect 4353 4573 4387 4607
rect 4905 4573 4939 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 7205 4573 7239 4607
rect 9137 4573 9171 4607
rect 10241 4573 10275 4607
rect 10334 4573 10368 4607
rect 10425 4573 10459 4607
rect 10977 4573 11011 4607
rect 11989 4573 12023 4607
rect 12081 4573 12115 4607
rect 12265 4573 12299 4607
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 14565 4573 14599 4607
rect 16129 4573 16163 4607
rect 16405 4573 16439 4607
rect 16865 4573 16899 4607
rect 17601 4573 17635 4607
rect 17785 4573 17819 4607
rect 18429 4573 18463 4607
rect 18705 4573 18739 4607
rect 19257 4573 19291 4607
rect 19350 4573 19384 4607
rect 19722 4573 19756 4607
rect 20545 4573 20579 4607
rect 8217 4505 8251 4539
rect 8401 4505 8435 4539
rect 11161 4505 11195 4539
rect 15301 4505 15335 4539
rect 16313 4505 16347 4539
rect 19533 4505 19567 4539
rect 19625 4505 19659 4539
rect 20729 4505 20763 4539
rect 2697 4437 2731 4471
rect 3985 4437 4019 4471
rect 4997 4437 5031 4471
rect 6377 4437 6411 4471
rect 7297 4437 7331 4471
rect 9413 4437 9447 4471
rect 14657 4437 14691 4471
rect 15393 4437 15427 4471
rect 18245 4437 18279 4471
rect 7021 4233 7055 4267
rect 8585 4233 8619 4267
rect 9505 4233 9539 4267
rect 9689 4233 9723 4267
rect 15945 4233 15979 4267
rect 17049 4233 17083 4267
rect 1869 4165 1903 4199
rect 2605 4165 2639 4199
rect 7757 4165 7791 4199
rect 10793 4165 10827 4199
rect 12081 4165 12115 4199
rect 12909 4165 12943 4199
rect 13737 4165 13771 4199
rect 17969 4165 18003 4199
rect 18153 4165 18187 4199
rect 19073 4165 19107 4199
rect 19901 4165 19935 4199
rect 3249 4097 3283 4131
rect 4060 4097 4094 4131
rect 4169 4097 4203 4131
rect 4445 4097 4479 4131
rect 4997 4097 5031 4131
rect 5641 4097 5675 4131
rect 6837 4097 6871 4131
rect 7113 4097 7147 4131
rect 8582 4097 8616 4131
rect 9686 4097 9720 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 11805 4097 11839 4131
rect 12633 4097 12667 4131
rect 12817 4097 12851 4131
rect 13001 4097 13035 4131
rect 14657 4097 14691 4131
rect 15669 4097 15703 4131
rect 15761 4097 15795 4131
rect 16037 4097 16071 4131
rect 16681 4097 16715 4131
rect 16773 4097 16807 4131
rect 18797 4097 18831 4131
rect 18981 4097 19015 4131
rect 19165 4097 19199 4131
rect 19809 4097 19843 4131
rect 20269 4097 20303 4131
rect 20545 4097 20579 4131
rect 2789 4029 2823 4063
rect 6653 4029 6687 4063
rect 9045 4029 9079 4063
rect 11621 4029 11655 4063
rect 12173 4029 12207 4063
rect 14841 4029 14875 4063
rect 18337 4029 18371 4063
rect 2053 3961 2087 3995
rect 3341 3961 3375 3995
rect 4353 3961 4387 3995
rect 5733 3961 5767 3995
rect 7941 3961 7975 3995
rect 13185 3961 13219 3995
rect 15577 3961 15611 3995
rect 20729 3961 20763 3995
rect 3893 3893 3927 3927
rect 5089 3893 5123 3927
rect 6377 3893 6411 3927
rect 6745 3893 6779 3927
rect 8401 3893 8435 3927
rect 8953 3893 8987 3927
rect 10885 3893 10919 3927
rect 11897 3893 11931 3927
rect 13829 3893 13863 3927
rect 15301 3893 15335 3927
rect 16773 3893 16807 3927
rect 19349 3893 19383 3927
rect 4445 3689 4479 3723
rect 6101 3689 6135 3723
rect 7205 3689 7239 3723
rect 9321 3689 9355 3723
rect 9873 3689 9907 3723
rect 10425 3689 10459 3723
rect 11713 3689 11747 3723
rect 12265 3689 12299 3723
rect 12909 3689 12943 3723
rect 14657 3689 14691 3723
rect 15669 3689 15703 3723
rect 18429 3689 18463 3723
rect 21649 4981 21683 5015
rect 21649 3893 21683 3927
rect 13461 3621 13495 3655
rect 17049 3621 17083 3655
rect 18337 3621 18371 3655
rect 20729 3621 20763 3655
rect 21557 3621 21591 3655
rect 5457 3553 5491 3587
rect 8217 3553 8251 3587
rect 11069 3553 11103 3587
rect 12357 3553 12391 3587
rect 17509 3553 17543 3587
rect 17693 3553 17727 3587
rect 18521 3553 18555 3587
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 6101 3485 6135 3519
rect 6285 3485 6319 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 9502 3485 9536 3519
rect 9965 3485 9999 3519
rect 10609 3485 10643 3519
rect 10701 3485 10735 3519
rect 11894 3485 11928 3519
rect 12817 3485 12851 3519
rect 13090 3485 13124 3519
rect 13553 3485 13587 3519
rect 14286 3485 14320 3519
rect 14749 3485 14783 3519
rect 15209 3485 15243 3519
rect 15393 3485 15427 3519
rect 15485 3485 15519 3519
rect 15761 3485 15795 3519
rect 18245 3485 18279 3519
rect 1869 3417 1903 3451
rect 3065 3417 3099 3451
rect 4169 3417 4203 3451
rect 5273 3417 5307 3451
rect 7757 3417 7791 3451
rect 10793 3417 10827 3451
rect 10911 3417 10945 3451
rect 16405 3417 16439 3451
rect 16589 3417 16623 3451
rect 19533 3417 19567 3451
rect 19809 3417 19843 3451
rect 19993 3417 20027 3451
rect 20545 3417 20579 3451
rect 1961 3349 1995 3383
rect 3157 3349 3191 3383
rect 4905 3349 4939 3383
rect 5365 3349 5399 3383
rect 6745 3349 6779 3383
rect 9505 3349 9539 3383
rect 11897 3349 11931 3383
rect 12817 3349 12851 3383
rect 13093 3349 13127 3383
rect 14105 3349 14139 3383
rect 14289 3349 14323 3383
rect 15209 3349 15243 3383
rect 17417 3349 17451 3383
rect 1501 3145 1535 3179
rect 4077 3145 4111 3179
rect 5273 3145 5307 3179
rect 5641 3145 5675 3179
rect 7021 3145 7055 3179
rect 8309 3145 8343 3179
rect 9597 3145 9631 3179
rect 10517 3145 10551 3179
rect 12081 3145 12115 3179
rect 14565 3145 14599 3179
rect 15669 3145 15703 3179
rect 15761 3145 15795 3179
rect 17969 3145 18003 3179
rect 18153 3145 18187 3179
rect 2237 3077 2271 3111
rect 3065 3077 3099 3111
rect 4169 3077 4203 3111
rect 7113 3077 7147 3111
rect 9229 3077 9263 3111
rect 10149 3077 10183 3111
rect 10333 3077 10367 3111
rect 12358 3077 12392 3111
rect 12567 3077 12601 3111
rect 13553 3077 13587 3111
rect 14473 3077 14507 3111
rect 16497 3077 16531 3111
rect 16773 3077 16807 3111
rect 20637 3077 20671 3111
rect 1685 3009 1719 3043
rect 3709 3009 3743 3043
rect 3893 3009 3927 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 8217 3009 8251 3043
rect 9045 3009 9079 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 12265 3009 12299 3043
rect 12449 3009 12483 3043
rect 12725 3009 12759 3043
rect 13185 3009 13219 3043
rect 13369 3009 13403 3043
rect 4261 2941 4295 2975
rect 7297 2941 7331 2975
rect 8401 2941 8435 2975
rect 14749 2941 14783 2975
rect 15853 2941 15887 2975
rect 3249 2873 3283 2907
rect 6653 2873 6687 2907
rect 15301 2873 15335 2907
rect 16497 2873 16531 2907
rect 16681 3009 16715 3043
rect 16957 3009 16991 3043
rect 18150 3009 18184 3043
rect 18521 3009 18555 3043
rect 19717 3009 19751 3043
rect 20453 3009 20487 3043
rect 17233 2941 17267 2975
rect 18613 2941 18647 2975
rect 2329 2805 2363 2839
rect 7849 2805 7883 2839
rect 14105 2805 14139 2839
rect 16681 2805 16715 2839
rect 17141 2805 17175 2839
rect 19809 2805 19843 2839
rect 5641 2601 5675 2635
rect 9505 2601 9539 2635
rect 16911 2601 16945 2635
rect 20637 2601 20671 2635
rect 2053 2533 2087 2567
rect 7021 2533 7055 2567
rect 15853 2533 15887 2567
rect 10425 2465 10459 2499
rect 12173 2465 12207 2499
rect 15117 2465 15151 2499
rect 18245 2465 18279 2499
rect 2789 2397 2823 2431
rect 5457 2397 5491 2431
rect 7757 2397 7791 2431
rect 10149 2397 10183 2431
rect 11897 2397 11931 2431
rect 14933 2397 14967 2431
rect 16681 2397 16715 2431
rect 19257 2397 19291 2431
rect 19533 2397 19567 2431
rect 20545 2397 20579 2431
rect 1869 2329 1903 2363
rect 2605 2329 2639 2363
rect 4261 2329 4295 2363
rect 6837 2329 6871 2363
rect 7573 2329 7607 2363
rect 9413 2329 9447 2363
rect 13277 2329 13311 2363
rect 15669 2329 15703 2363
rect 18061 2329 18095 2363
rect 4353 2261 4387 2295
rect 13369 2261 13403 2295
<< metal1 >>
rect 17862 22448 17868 22500
rect 17920 22488 17926 22500
rect 18322 22488 18328 22500
rect 17920 22460 18328 22488
rect 17920 22448 17926 22460
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 1104 22330 21436 22352
rect 1104 22278 4338 22330
rect 4390 22278 4402 22330
rect 4454 22278 4466 22330
rect 4518 22278 4530 22330
rect 4582 22278 4594 22330
rect 4646 22278 11116 22330
rect 11168 22278 11180 22330
rect 11232 22278 11244 22330
rect 11296 22278 11308 22330
rect 11360 22278 11372 22330
rect 11424 22278 17893 22330
rect 17945 22278 17957 22330
rect 18009 22278 18021 22330
rect 18073 22278 18085 22330
rect 18137 22278 18149 22330
rect 18201 22278 21436 22330
rect 1104 22256 21436 22278
rect 14826 22216 14832 22228
rect 14660 22188 14832 22216
rect 5350 22108 5356 22160
rect 5408 22148 5414 22160
rect 6365 22151 6423 22157
rect 6365 22148 6377 22151
rect 5408 22120 6377 22148
rect 5408 22108 5414 22120
rect 6365 22117 6377 22120
rect 6411 22117 6423 22151
rect 6365 22111 6423 22117
rect 4062 22040 4068 22092
rect 4120 22080 4126 22092
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 4120 22052 4169 22080
rect 4120 22040 4126 22052
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 5718 22040 5724 22092
rect 5776 22080 5782 22092
rect 6825 22083 6883 22089
rect 6825 22080 6837 22083
rect 5776 22052 6837 22080
rect 5776 22040 5782 22052
rect 6825 22049 6837 22052
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 7929 22083 7987 22089
rect 7929 22049 7941 22083
rect 7975 22080 7987 22083
rect 7975 22052 11100 22080
rect 7975 22049 7987 22052
rect 7929 22043 7987 22049
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2774 22012 2780 22024
rect 1903 21984 2780 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3510 22012 3516 22024
rect 3099 21984 3516 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 3510 21972 3516 21984
rect 3568 21972 3574 22024
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 21981 4491 22015
rect 4433 21975 4491 21981
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 22012 5687 22015
rect 5902 22012 5908 22024
rect 5675 21984 5908 22012
rect 5675 21981 5687 21984
rect 5629 21975 5687 21981
rect 3237 21947 3295 21953
rect 3237 21913 3249 21947
rect 3283 21944 3295 21947
rect 3602 21944 3608 21956
rect 3283 21916 3608 21944
rect 3283 21913 3295 21916
rect 3237 21907 3295 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 4448 21944 4476 21975
rect 5902 21972 5908 21984
rect 5960 21972 5966 22024
rect 6270 21972 6276 22024
rect 6328 22012 6334 22024
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 6328 21984 6561 22012
rect 6328 21972 6334 21984
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 6914 22012 6920 22024
rect 6696 21984 6741 22012
rect 6875 21984 6920 22012
rect 6696 21972 6702 21984
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 7616 21984 7757 22012
rect 7616 21972 7622 21984
rect 7745 21981 7757 21984
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 8352 21984 9413 22012
rect 8352 21972 8358 21984
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 10008 21984 10057 22012
rect 10008 21972 10014 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10781 22015 10839 22021
rect 10781 22012 10793 22015
rect 10652 21984 10793 22012
rect 10652 21972 10658 21984
rect 10781 21981 10793 21984
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 10870 21972 10876 22024
rect 10928 22012 10934 22024
rect 10965 22015 11023 22021
rect 10965 22012 10977 22015
rect 10928 21984 10977 22012
rect 10928 21972 10934 21984
rect 10965 21981 10977 21984
rect 11011 21981 11023 22015
rect 11072 22012 11100 22052
rect 11146 22040 11152 22092
rect 11204 22080 11210 22092
rect 11517 22083 11575 22089
rect 11517 22080 11529 22083
rect 11204 22052 11529 22080
rect 11204 22040 11210 22052
rect 11517 22049 11529 22052
rect 11563 22049 11575 22083
rect 14660 22080 14688 22188
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 11517 22043 11575 22049
rect 11624 22052 14688 22080
rect 11624 22012 11652 22052
rect 14734 22040 14740 22092
rect 14792 22080 14798 22092
rect 14829 22083 14887 22089
rect 14829 22080 14841 22083
rect 14792 22052 14841 22080
rect 14792 22040 14798 22052
rect 14829 22049 14841 22052
rect 14875 22049 14887 22083
rect 15378 22080 15384 22092
rect 14829 22043 14887 22049
rect 15028 22052 15384 22080
rect 11072 21984 11652 22012
rect 10965 21975 11023 21981
rect 11698 21972 11704 22024
rect 11756 22012 11762 22024
rect 11793 22015 11851 22021
rect 11793 22012 11805 22015
rect 11756 21984 11805 22012
rect 11756 21972 11762 21984
rect 11793 21981 11805 21984
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12897 22015 12955 22021
rect 12897 22012 12909 22015
rect 12492 21984 12909 22012
rect 12492 21972 12498 21984
rect 12897 21981 12909 21984
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 22012 14243 22015
rect 15028 22012 15056 22052
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17313 22083 17371 22089
rect 17313 22080 17325 22083
rect 16908 22052 17325 22080
rect 16908 22040 16914 22052
rect 17313 22049 17325 22052
rect 17359 22049 17371 22083
rect 17313 22043 17371 22049
rect 17402 22040 17408 22092
rect 17460 22080 17466 22092
rect 19889 22083 19947 22089
rect 17460 22052 19472 22080
rect 17460 22040 17466 22052
rect 14231 21984 15056 22012
rect 14231 21981 14243 21984
rect 14185 21975 14243 21981
rect 15102 21972 15108 22024
rect 15160 22012 15166 22024
rect 15160 21984 15205 22012
rect 15160 21972 15166 21984
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 17129 22015 17187 22021
rect 17129 22012 17141 22015
rect 16632 21984 17141 22012
rect 16632 21972 16638 21984
rect 17129 21981 17141 21984
rect 17175 21981 17187 22015
rect 18506 22012 18512 22024
rect 18467 21984 18512 22012
rect 17129 21975 17187 21981
rect 18506 21972 18512 21984
rect 18564 21972 18570 22024
rect 19444 22021 19472 22052
rect 19889 22049 19901 22083
rect 19935 22080 19947 22083
rect 21358 22080 21364 22092
rect 19935 22052 21364 22080
rect 19935 22049 19947 22052
rect 19889 22043 19947 22049
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 20162 22012 20168 22024
rect 20123 21984 20168 22012
rect 19429 21975 19487 21981
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 14369 21947 14427 21953
rect 4448 21916 6500 21944
rect 1949 21879 2007 21885
rect 1949 21845 1961 21879
rect 1995 21876 2007 21879
rect 5534 21876 5540 21888
rect 1995 21848 5540 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 5721 21879 5779 21885
rect 5721 21845 5733 21879
rect 5767 21876 5779 21879
rect 5994 21876 6000 21888
rect 5767 21848 6000 21876
rect 5767 21845 5779 21848
rect 5721 21839 5779 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6472 21876 6500 21916
rect 8404 21916 14136 21944
rect 8404 21876 8432 21916
rect 6472 21848 8432 21876
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 9493 21879 9551 21885
rect 9493 21876 9505 21879
rect 8996 21848 9505 21876
rect 8996 21836 9002 21848
rect 9493 21845 9505 21848
rect 9539 21845 9551 21879
rect 9493 21839 9551 21845
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 10502 21876 10508 21888
rect 10275 21848 10508 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10870 21876 10876 21888
rect 10831 21848 10876 21876
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 12216 21848 13001 21876
rect 12216 21836 12222 21848
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 14108 21876 14136 21916
rect 14369 21913 14381 21947
rect 14415 21944 14427 21947
rect 18966 21944 18972 21956
rect 14415 21916 18972 21944
rect 14415 21913 14427 21916
rect 14369 21907 14427 21913
rect 18966 21904 18972 21916
rect 19024 21904 19030 21956
rect 17034 21876 17040 21888
rect 14108 21848 17040 21876
rect 12989 21839 13047 21845
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17218 21836 17224 21888
rect 17276 21876 17282 21888
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 17276 21848 18613 21876
rect 17276 21836 17282 21848
rect 18601 21845 18613 21848
rect 18647 21845 18659 21879
rect 18601 21839 18659 21845
rect 19245 21879 19303 21885
rect 19245 21845 19257 21879
rect 19291 21876 19303 21879
rect 19334 21876 19340 21888
rect 19291 21848 19340 21876
rect 19291 21845 19303 21848
rect 19245 21839 19303 21845
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 1104 21786 21436 21808
rect 1104 21734 7727 21786
rect 7779 21734 7791 21786
rect 7843 21734 7855 21786
rect 7907 21734 7919 21786
rect 7971 21734 7983 21786
rect 8035 21734 14504 21786
rect 14556 21734 14568 21786
rect 14620 21734 14632 21786
rect 14684 21734 14696 21786
rect 14748 21734 14760 21786
rect 14812 21734 21436 21786
rect 1104 21712 21436 21734
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4295 21644 4997 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 4985 21641 4997 21644
rect 5031 21641 5043 21675
rect 4985 21635 5043 21641
rect 5169 21675 5227 21681
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5350 21672 5356 21684
rect 5215 21644 5356 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 6733 21675 6791 21681
rect 6733 21641 6745 21675
rect 6779 21672 6791 21675
rect 8389 21675 8447 21681
rect 8389 21672 8401 21675
rect 6779 21644 8401 21672
rect 6779 21641 6791 21644
rect 6733 21635 6791 21641
rect 8389 21641 8401 21644
rect 8435 21641 8447 21675
rect 8389 21635 8447 21641
rect 9398 21632 9404 21684
rect 9456 21672 9462 21684
rect 9493 21675 9551 21681
rect 9493 21672 9505 21675
rect 9456 21644 9505 21672
rect 9456 21632 9462 21644
rect 9493 21641 9505 21644
rect 9539 21641 9551 21675
rect 10226 21672 10232 21684
rect 9493 21635 9551 21641
rect 9646 21644 10232 21672
rect 1854 21604 1860 21616
rect 1815 21576 1860 21604
rect 1854 21564 1860 21576
rect 1912 21564 1918 21616
rect 2041 21607 2099 21613
rect 2041 21573 2053 21607
rect 2087 21604 2099 21607
rect 4890 21604 4896 21616
rect 2087 21576 4896 21604
rect 2087 21573 2099 21576
rect 2041 21567 2099 21573
rect 4890 21564 4896 21576
rect 4948 21564 4954 21616
rect 6825 21607 6883 21613
rect 6825 21604 6837 21607
rect 6564 21576 6837 21604
rect 6564 21548 6592 21576
rect 6825 21573 6837 21576
rect 6871 21573 6883 21607
rect 6825 21567 6883 21573
rect 9306 21564 9312 21616
rect 9364 21604 9370 21616
rect 9646 21604 9674 21644
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11572 21644 11713 21672
rect 11572 21632 11578 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 12437 21675 12495 21681
rect 12437 21641 12449 21675
rect 12483 21672 12495 21675
rect 13722 21672 13728 21684
rect 12483 21644 13728 21672
rect 12483 21641 12495 21644
rect 12437 21635 12495 21641
rect 9364 21576 9674 21604
rect 9364 21564 9370 21576
rect 11422 21564 11428 21616
rect 11480 21604 11486 21616
rect 12452 21604 12480 21635
rect 13722 21632 13728 21644
rect 13780 21672 13786 21684
rect 13780 21644 14412 21672
rect 13780 21632 13786 21644
rect 13078 21604 13084 21616
rect 11480 21576 12480 21604
rect 12544 21576 13084 21604
rect 11480 21564 11486 21576
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 3142 21536 3148 21548
rect 2547 21508 3148 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 4157 21539 4215 21545
rect 4157 21505 4169 21539
rect 4203 21505 4215 21539
rect 4157 21499 4215 21505
rect 5166 21539 5224 21545
rect 5166 21505 5178 21539
rect 5212 21536 5224 21539
rect 5442 21536 5448 21548
rect 5212 21508 5448 21536
rect 5212 21505 5224 21508
rect 5166 21499 5224 21505
rect 1762 21360 1768 21412
rect 1820 21400 1826 21412
rect 2685 21403 2743 21409
rect 2685 21400 2697 21403
rect 1820 21372 2697 21400
rect 1820 21360 1826 21372
rect 2685 21369 2697 21372
rect 2731 21369 2743 21403
rect 2685 21363 2743 21369
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3108 21304 3801 21332
rect 3108 21292 3114 21304
rect 3789 21301 3801 21304
rect 3835 21301 3847 21335
rect 4172 21332 4200 21499
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 6178 21536 6184 21548
rect 5675 21508 6184 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 6546 21536 6552 21548
rect 6507 21508 6552 21536
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 8294 21536 8300 21548
rect 8255 21508 8300 21536
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21536 9459 21539
rect 10042 21536 10048 21548
rect 9447 21508 10048 21536
rect 9447 21505 9459 21508
rect 9401 21499 9459 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10226 21496 10232 21548
rect 10284 21536 10290 21548
rect 11609 21539 11667 21545
rect 10284 21508 10329 21536
rect 10284 21496 10290 21508
rect 11609 21505 11621 21539
rect 11655 21505 11667 21539
rect 11609 21499 11667 21505
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 12342 21536 12348 21548
rect 12299 21508 12348 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 4433 21471 4491 21477
rect 4433 21437 4445 21471
rect 4479 21437 4491 21471
rect 4433 21431 4491 21437
rect 4448 21400 4476 21431
rect 5350 21428 5356 21480
rect 5408 21468 5414 21480
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 5408 21440 5549 21468
rect 5408 21428 5414 21440
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 5644 21440 6316 21468
rect 5644 21400 5672 21440
rect 4448 21372 5672 21400
rect 6288 21400 6316 21440
rect 6362 21428 6368 21480
rect 6420 21468 6426 21480
rect 6917 21471 6975 21477
rect 6917 21468 6929 21471
rect 6420 21440 6929 21468
rect 6420 21428 6426 21440
rect 6917 21437 6929 21440
rect 6963 21437 6975 21471
rect 7466 21468 7472 21480
rect 6917 21431 6975 21437
rect 7024 21440 7472 21468
rect 7024 21400 7052 21440
rect 7466 21428 7472 21440
rect 7524 21468 7530 21480
rect 8018 21468 8024 21480
rect 7524 21440 8024 21468
rect 7524 21428 7530 21440
rect 8018 21428 8024 21440
rect 8076 21468 8082 21480
rect 8481 21471 8539 21477
rect 8481 21468 8493 21471
rect 8076 21440 8493 21468
rect 8076 21428 8082 21440
rect 8481 21437 8493 21440
rect 8527 21468 8539 21471
rect 8527 21440 8800 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 6288 21372 7052 21400
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 7929 21403 7987 21409
rect 7929 21400 7941 21403
rect 7616 21372 7941 21400
rect 7616 21360 7622 21372
rect 7929 21369 7941 21372
rect 7975 21369 7987 21403
rect 7929 21363 7987 21369
rect 8662 21332 8668 21344
rect 4172 21304 8668 21332
rect 3789 21295 3847 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8772 21332 8800 21440
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 9272 21440 10517 21468
rect 9272 21428 9278 21440
rect 10505 21437 10517 21440
rect 10551 21468 10563 21471
rect 11514 21468 11520 21480
rect 10551 21440 11520 21468
rect 10551 21437 10563 21440
rect 10505 21431 10563 21437
rect 11514 21428 11520 21440
rect 11572 21428 11578 21480
rect 11624 21468 11652 21499
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 12544 21545 12572 21576
rect 13078 21564 13084 21576
rect 13136 21604 13142 21616
rect 13262 21604 13268 21616
rect 13136 21576 13268 21604
rect 13136 21564 13142 21576
rect 13262 21564 13268 21576
rect 13320 21564 13326 21616
rect 13357 21607 13415 21613
rect 13357 21573 13369 21607
rect 13403 21573 13415 21607
rect 13357 21567 13415 21573
rect 12529 21539 12587 21545
rect 12529 21505 12541 21539
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 13170 21496 13176 21548
rect 13228 21536 13234 21548
rect 13372 21536 13400 21567
rect 13446 21564 13452 21616
rect 13504 21604 13510 21616
rect 13504 21576 14228 21604
rect 13504 21564 13510 21576
rect 13814 21536 13820 21548
rect 13228 21508 13400 21536
rect 13556 21508 13820 21536
rect 13228 21496 13234 21508
rect 13262 21468 13268 21480
rect 11624 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 13446 21468 13452 21480
rect 13407 21440 13452 21468
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 13556 21477 13584 21508
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14200 21545 14228 21576
rect 14384 21545 14412 21644
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 14884 21644 16988 21672
rect 14884 21632 14890 21644
rect 14458 21564 14464 21616
rect 14516 21604 14522 21616
rect 15933 21607 15991 21613
rect 15933 21604 15945 21607
rect 14516 21576 15945 21604
rect 14516 21564 14522 21576
rect 15933 21573 15945 21576
rect 15979 21573 15991 21607
rect 15933 21567 15991 21573
rect 16022 21564 16028 21616
rect 16080 21604 16086 21616
rect 16853 21607 16911 21613
rect 16853 21604 16865 21607
rect 16080 21576 16865 21604
rect 16080 21564 16086 21576
rect 16853 21573 16865 21576
rect 16899 21573 16911 21607
rect 16960 21604 16988 21644
rect 17034 21632 17040 21684
rect 17092 21672 17098 21684
rect 17865 21675 17923 21681
rect 17865 21672 17877 21675
rect 17092 21644 17877 21672
rect 17092 21632 17098 21644
rect 17865 21641 17877 21644
rect 17911 21672 17923 21675
rect 17911 21644 18644 21672
rect 17911 21641 17923 21644
rect 17865 21635 17923 21641
rect 18616 21613 18644 21644
rect 18601 21607 18659 21613
rect 16960 21576 18552 21604
rect 16853 21567 16911 21573
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21505 14243 21539
rect 14185 21499 14243 21505
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21505 14887 21539
rect 15010 21536 15016 21548
rect 14971 21508 15016 21536
rect 14829 21499 14887 21505
rect 13541 21471 13599 21477
rect 13541 21437 13553 21471
rect 13587 21437 13599 21471
rect 13541 21431 13599 21437
rect 13630 21428 13636 21480
rect 13688 21468 13694 21480
rect 14844 21468 14872 21499
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 15838 21536 15844 21548
rect 15243 21508 15844 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 13688 21440 14872 21468
rect 15120 21468 15148 21499
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 17494 21496 17500 21548
rect 17552 21536 17558 21548
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17552 21508 17693 21536
rect 17552 21496 17558 21508
rect 17681 21505 17693 21508
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21536 18015 21539
rect 18230 21536 18236 21548
rect 18003 21508 18236 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 18230 21496 18236 21508
rect 18288 21536 18294 21548
rect 18417 21539 18475 21545
rect 18417 21536 18429 21539
rect 18288 21508 18429 21536
rect 18288 21496 18294 21508
rect 18417 21505 18429 21508
rect 18463 21505 18475 21539
rect 18524 21536 18552 21576
rect 18601 21573 18613 21607
rect 18647 21604 18659 21607
rect 18647 21576 19288 21604
rect 18647 21573 18659 21576
rect 18601 21567 18659 21573
rect 19058 21536 19064 21548
rect 18524 21508 19064 21536
rect 18417 21499 18475 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19260 21545 19288 21576
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21505 19303 21539
rect 19245 21499 19303 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 22462 21536 22468 21548
rect 19935 21508 22468 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 15286 21468 15292 21480
rect 15120 21440 15292 21468
rect 13688 21428 13694 21440
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 16117 21471 16175 21477
rect 16117 21468 16129 21471
rect 15528 21440 16129 21468
rect 15528 21428 15534 21440
rect 16117 21437 16129 21440
rect 16163 21437 16175 21471
rect 16117 21431 16175 21437
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 20165 21471 20223 21477
rect 20165 21468 20177 21471
rect 19484 21440 20177 21468
rect 19484 21428 19490 21440
rect 20165 21437 20177 21440
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 9122 21360 9128 21412
rect 9180 21400 9186 21412
rect 12989 21403 13047 21409
rect 12989 21400 13001 21403
rect 9180 21372 13001 21400
rect 9180 21360 9186 21372
rect 12989 21369 13001 21372
rect 13035 21369 13047 21403
rect 12989 21363 13047 21369
rect 13170 21360 13176 21412
rect 13228 21400 13234 21412
rect 16574 21400 16580 21412
rect 13228 21372 16580 21400
rect 13228 21360 13234 21372
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 17037 21403 17095 21409
rect 17037 21369 17049 21403
rect 17083 21400 17095 21403
rect 17402 21400 17408 21412
rect 17083 21372 17408 21400
rect 17083 21369 17095 21372
rect 17037 21363 17095 21369
rect 17402 21360 17408 21372
rect 17460 21360 17466 21412
rect 17586 21360 17592 21412
rect 17644 21400 17650 21412
rect 19337 21403 19395 21409
rect 19337 21400 19349 21403
rect 17644 21372 19349 21400
rect 17644 21360 17650 21372
rect 19337 21369 19349 21372
rect 19383 21369 19395 21403
rect 19337 21363 19395 21369
rect 9950 21332 9956 21344
rect 8772 21304 9956 21332
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10045 21335 10103 21341
rect 10045 21301 10057 21335
rect 10091 21332 10103 21335
rect 10318 21332 10324 21344
rect 10091 21304 10324 21332
rect 10091 21301 10103 21304
rect 10045 21295 10103 21301
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 10410 21292 10416 21344
rect 10468 21332 10474 21344
rect 10468 21304 10513 21332
rect 10468 21292 10474 21304
rect 11514 21292 11520 21344
rect 11572 21332 11578 21344
rect 11974 21332 11980 21344
rect 11572 21304 11980 21332
rect 11572 21292 11578 21304
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 12250 21332 12256 21344
rect 12211 21304 12256 21332
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12342 21292 12348 21344
rect 12400 21332 12406 21344
rect 12894 21332 12900 21344
rect 12400 21304 12900 21332
rect 12400 21292 12406 21304
rect 12894 21292 12900 21304
rect 12952 21332 12958 21344
rect 14185 21335 14243 21341
rect 14185 21332 14197 21335
rect 12952 21304 14197 21332
rect 12952 21292 12958 21304
rect 14185 21301 14197 21304
rect 14231 21301 14243 21335
rect 14185 21295 14243 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15381 21335 15439 21341
rect 15381 21332 15393 21335
rect 15068 21304 15393 21332
rect 15068 21292 15074 21304
rect 15381 21301 15393 21304
rect 15427 21301 15439 21335
rect 15381 21295 15439 21301
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 17218 21332 17224 21344
rect 15528 21304 17224 21332
rect 15528 21292 15534 21304
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 17497 21335 17555 21341
rect 17497 21301 17509 21335
rect 17543 21332 17555 21335
rect 17770 21332 17776 21344
rect 17543 21304 17776 21332
rect 17543 21301 17555 21304
rect 17497 21295 17555 21301
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 18506 21292 18512 21344
rect 18564 21332 18570 21344
rect 18785 21335 18843 21341
rect 18785 21332 18797 21335
rect 18564 21304 18797 21332
rect 18564 21292 18570 21304
rect 18785 21301 18797 21304
rect 18831 21301 18843 21335
rect 18785 21295 18843 21301
rect 1104 21242 21436 21264
rect 1104 21190 4338 21242
rect 4390 21190 4402 21242
rect 4454 21190 4466 21242
rect 4518 21190 4530 21242
rect 4582 21190 4594 21242
rect 4646 21190 11116 21242
rect 11168 21190 11180 21242
rect 11232 21190 11244 21242
rect 11296 21190 11308 21242
rect 11360 21190 11372 21242
rect 11424 21190 17893 21242
rect 17945 21190 17957 21242
rect 18009 21190 18021 21242
rect 18073 21190 18085 21242
rect 18137 21190 18149 21242
rect 18201 21190 21436 21242
rect 1104 21168 21436 21190
rect 566 21088 572 21140
rect 624 21128 630 21140
rect 1949 21131 2007 21137
rect 1949 21128 1961 21131
rect 624 21100 1961 21128
rect 624 21088 630 21100
rect 1949 21097 1961 21100
rect 1995 21097 2007 21131
rect 1949 21091 2007 21097
rect 4706 21088 4712 21140
rect 4764 21128 4770 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 4764 21100 6929 21128
rect 4764 21088 4770 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21128 7987 21131
rect 8018 21128 8024 21140
rect 7975 21100 8024 21128
rect 7975 21097 7987 21100
rect 7929 21091 7987 21097
rect 8018 21088 8024 21100
rect 8076 21088 8082 21140
rect 9309 21131 9367 21137
rect 9309 21097 9321 21131
rect 9355 21128 9367 21131
rect 9858 21128 9864 21140
rect 9355 21100 9864 21128
rect 9355 21097 9367 21100
rect 9309 21091 9367 21097
rect 9858 21088 9864 21100
rect 9916 21128 9922 21140
rect 10870 21128 10876 21140
rect 9916 21100 10876 21128
rect 9916 21088 9922 21100
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 11606 21088 11612 21140
rect 11664 21128 11670 21140
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11664 21100 11713 21128
rect 11664 21088 11670 21100
rect 11701 21097 11713 21100
rect 11747 21097 11759 21131
rect 11701 21091 11759 21097
rect 12897 21131 12955 21137
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 13354 21128 13360 21140
rect 12943 21100 13360 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 13449 21131 13507 21137
rect 13449 21097 13461 21131
rect 13495 21128 13507 21131
rect 13630 21128 13636 21140
rect 13495 21100 13636 21128
rect 13495 21097 13507 21100
rect 13449 21091 13507 21097
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 14366 21128 14372 21140
rect 14327 21100 14372 21128
rect 14366 21088 14372 21100
rect 14424 21088 14430 21140
rect 16390 21128 16396 21140
rect 16351 21100 16396 21128
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 2222 21020 2228 21072
rect 2280 21060 2286 21072
rect 2777 21063 2835 21069
rect 2777 21060 2789 21063
rect 2280 21032 2789 21060
rect 2280 21020 2286 21032
rect 2777 21029 2789 21032
rect 2823 21029 2835 21063
rect 2777 21023 2835 21029
rect 3789 21063 3847 21069
rect 3789 21029 3801 21063
rect 3835 21060 3847 21063
rect 4982 21060 4988 21072
rect 3835 21032 4988 21060
rect 3835 21029 3847 21032
rect 3789 21023 3847 21029
rect 4982 21020 4988 21032
rect 5040 21060 5046 21072
rect 5040 21032 6156 21060
rect 5040 21020 5046 21032
rect 4338 20992 4344 21004
rect 4299 20964 4344 20992
rect 4338 20952 4344 20964
rect 4396 20952 4402 21004
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 5868 20964 6040 20992
rect 5868 20952 5874 20964
rect 1118 20884 1124 20936
rect 1176 20924 1182 20936
rect 5261 20927 5319 20933
rect 5261 20924 5273 20927
rect 1176 20896 5273 20924
rect 1176 20884 1182 20896
rect 5261 20893 5273 20896
rect 5307 20893 5319 20927
rect 5261 20887 5319 20893
rect 5534 20884 5540 20936
rect 5592 20884 5598 20936
rect 5718 20924 5724 20936
rect 5679 20896 5724 20924
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 5902 20924 5908 20936
rect 5863 20896 5908 20924
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 6012 20933 6040 20964
rect 6128 20933 6156 21032
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 7837 21063 7895 21069
rect 7837 21060 7849 21063
rect 7248 21032 7849 21060
rect 7248 21020 7254 21032
rect 7837 21029 7849 21032
rect 7883 21060 7895 21063
rect 9953 21063 10011 21069
rect 7883 21032 9720 21060
rect 7883 21029 7895 21032
rect 7837 21023 7895 21029
rect 8478 20992 8484 21004
rect 8036 20964 8484 20992
rect 8036 20933 8064 20964
rect 8478 20952 8484 20964
rect 8536 20992 8542 21004
rect 9493 20995 9551 21001
rect 8536 20964 9352 20992
rect 8536 20952 8542 20964
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 6128 20927 6193 20933
rect 6128 20896 6147 20927
rect 5997 20887 6055 20893
rect 6135 20893 6147 20896
rect 6181 20893 6193 20927
rect 6135 20887 6193 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7745 20927 7803 20933
rect 6871 20896 7696 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 1857 20859 1915 20865
rect 1857 20825 1869 20859
rect 1903 20856 1915 20859
rect 2498 20856 2504 20868
rect 1903 20828 2504 20856
rect 1903 20825 1915 20828
rect 1857 20819 1915 20825
rect 2498 20816 2504 20828
rect 2556 20816 2562 20868
rect 2593 20859 2651 20865
rect 2593 20825 2605 20859
rect 2639 20856 2651 20859
rect 2639 20828 5028 20856
rect 2639 20825 2651 20828
rect 2593 20819 2651 20825
rect 4154 20788 4160 20800
rect 4115 20760 4160 20788
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 4246 20748 4252 20800
rect 4304 20788 4310 20800
rect 5000 20788 5028 20828
rect 5074 20816 5080 20868
rect 5132 20856 5138 20868
rect 5552 20856 5580 20884
rect 6362 20856 6368 20868
rect 5132 20828 5177 20856
rect 5552 20828 6368 20856
rect 5132 20816 5138 20828
rect 6362 20816 6368 20828
rect 6420 20816 6426 20868
rect 7668 20856 7696 20896
rect 7745 20893 7757 20927
rect 7791 20924 7803 20927
rect 8021 20927 8079 20933
rect 7791 20896 7880 20924
rect 7791 20893 7803 20896
rect 7745 20887 7803 20893
rect 7852 20856 7880 20896
rect 8021 20893 8033 20927
rect 8067 20893 8079 20927
rect 8202 20924 8208 20936
rect 8163 20896 8208 20924
rect 8021 20887 8079 20893
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 9214 20924 9220 20936
rect 9175 20896 9220 20924
rect 9214 20884 9220 20896
rect 9272 20884 9278 20936
rect 8110 20856 8116 20868
rect 7668 20828 7788 20856
rect 7852 20828 8116 20856
rect 5534 20788 5540 20800
rect 4304 20760 4349 20788
rect 5000 20760 5540 20788
rect 4304 20748 4310 20760
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 5626 20748 5632 20800
rect 5684 20788 5690 20800
rect 6270 20788 6276 20800
rect 5684 20760 6276 20788
rect 5684 20748 5690 20760
rect 6270 20748 6276 20760
rect 6328 20748 6334 20800
rect 7469 20791 7527 20797
rect 7469 20757 7481 20791
rect 7515 20788 7527 20791
rect 7650 20788 7656 20800
rect 7515 20760 7656 20788
rect 7515 20757 7527 20760
rect 7469 20751 7527 20757
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 7760 20788 7788 20828
rect 8110 20816 8116 20828
rect 8168 20816 8174 20868
rect 9122 20788 9128 20800
rect 7760 20760 9128 20788
rect 9122 20748 9128 20760
rect 9180 20748 9186 20800
rect 9324 20788 9352 20964
rect 9493 20961 9505 20995
rect 9539 20992 9551 20995
rect 9582 20992 9588 21004
rect 9539 20964 9588 20992
rect 9539 20961 9551 20964
rect 9493 20955 9551 20961
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9692 20924 9720 21032
rect 9953 21029 9965 21063
rect 9999 21060 10011 21063
rect 11885 21063 11943 21069
rect 9999 21032 11008 21060
rect 9999 21029 10011 21032
rect 9953 21023 10011 21029
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 10410 20992 10416 21004
rect 9824 20964 10416 20992
rect 9824 20952 9830 20964
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 10597 20995 10655 21001
rect 10597 20961 10609 20995
rect 10643 20992 10655 20995
rect 10778 20992 10784 21004
rect 10643 20964 10784 20992
rect 10643 20961 10655 20964
rect 10597 20955 10655 20961
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 10134 20924 10140 20936
rect 9692 20896 10140 20924
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 10376 20896 10421 20924
rect 10376 20884 10382 20896
rect 9493 20859 9551 20865
rect 9493 20825 9505 20859
rect 9539 20856 9551 20859
rect 10980 20856 11008 21032
rect 11885 21029 11897 21063
rect 11931 21029 11943 21063
rect 11885 21023 11943 21029
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11793 20995 11851 21001
rect 11793 20992 11805 20995
rect 11112 20964 11805 20992
rect 11112 20952 11118 20964
rect 11793 20961 11805 20964
rect 11839 20961 11851 20995
rect 11900 20992 11928 21023
rect 15838 21020 15844 21072
rect 15896 21060 15902 21072
rect 17313 21063 17371 21069
rect 17313 21060 17325 21063
rect 15896 21032 17325 21060
rect 15896 21020 15902 21032
rect 17313 21029 17325 21032
rect 17359 21029 17371 21063
rect 17313 21023 17371 21029
rect 12526 20992 12532 21004
rect 11900 20964 12532 20992
rect 11793 20955 11851 20961
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 15013 20995 15071 21001
rect 15013 20992 15025 20995
rect 13872 20964 15025 20992
rect 13872 20952 13878 20964
rect 15013 20961 15025 20964
rect 15059 20992 15071 20995
rect 15059 20964 15516 20992
rect 15059 20961 15071 20964
rect 15013 20955 15071 20961
rect 11974 20884 11980 20936
rect 12032 20924 12038 20936
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 12032 20896 12173 20924
rect 12032 20884 12038 20896
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 13078 20927 13136 20933
rect 13078 20893 13090 20927
rect 13124 20924 13136 20927
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13124 20896 13553 20924
rect 13124 20893 13136 20896
rect 13078 20887 13136 20893
rect 13541 20893 13553 20896
rect 13587 20924 13599 20927
rect 13998 20924 14004 20936
rect 13587 20896 14004 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 13998 20884 14004 20896
rect 14056 20924 14062 20936
rect 15102 20924 15108 20936
rect 14056 20896 15108 20924
rect 14056 20884 14062 20896
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 15488 20924 15516 20964
rect 16114 20952 16120 21004
rect 16172 20992 16178 21004
rect 16485 20995 16543 21001
rect 16485 20992 16497 20995
rect 16172 20964 16497 20992
rect 16172 20952 16178 20964
rect 16485 20961 16497 20964
rect 16531 20961 16543 20995
rect 16485 20955 16543 20961
rect 16577 20995 16635 21001
rect 16577 20961 16589 20995
rect 16623 20992 16635 20995
rect 16942 20992 16948 21004
rect 16623 20964 16948 20992
rect 16623 20961 16635 20964
rect 16577 20955 16635 20961
rect 16592 20924 16620 20955
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 17770 20992 17776 21004
rect 17731 20964 17776 20992
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 17920 20964 17965 20992
rect 17920 20952 17926 20964
rect 15488 20896 16620 20924
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20924 16727 20927
rect 16758 20924 16764 20936
rect 16715 20896 16764 20924
rect 16715 20893 16727 20896
rect 16669 20887 16727 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20924 16911 20927
rect 17586 20924 17592 20936
rect 16899 20896 17592 20924
rect 16899 20893 16911 20896
rect 16853 20887 16911 20893
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 18506 20924 18512 20936
rect 18467 20896 18512 20924
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 19518 20884 19524 20936
rect 19576 20924 19582 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19576 20896 19625 20924
rect 19576 20884 19582 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 21910 20924 21916 20936
rect 20487 20896 21916 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 21910 20884 21916 20896
rect 21968 20884 21974 20936
rect 13170 20856 13176 20868
rect 9539 20828 10180 20856
rect 10980 20828 13176 20856
rect 9539 20825 9551 20828
rect 9493 20819 9551 20825
rect 10152 20822 10180 20828
rect 10042 20788 10048 20800
rect 9324 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10152 20797 10456 20822
rect 13170 20816 13176 20828
rect 13228 20816 13234 20868
rect 13262 20816 13268 20868
rect 13320 20856 13326 20868
rect 13446 20856 13452 20868
rect 13320 20828 13452 20856
rect 13320 20816 13326 20828
rect 13446 20816 13452 20828
rect 13504 20816 13510 20868
rect 14458 20816 14464 20868
rect 14516 20816 14522 20868
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 15562 20856 15568 20868
rect 14783 20828 15568 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 17494 20816 17500 20868
rect 17552 20856 17558 20868
rect 18601 20859 18659 20865
rect 18601 20856 18613 20859
rect 17552 20828 18613 20856
rect 17552 20816 17558 20828
rect 18601 20825 18613 20828
rect 18647 20825 18659 20859
rect 18601 20819 18659 20825
rect 10152 20794 10471 20797
rect 10413 20791 10471 20794
rect 10413 20757 10425 20791
rect 10459 20757 10471 20791
rect 10413 20751 10471 20757
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11606 20788 11612 20800
rect 11471 20760 11612 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 12066 20788 12072 20800
rect 12027 20760 12072 20788
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 13081 20791 13139 20797
rect 13081 20788 13093 20791
rect 12492 20760 13093 20788
rect 12492 20748 12498 20760
rect 13081 20757 13093 20760
rect 13127 20788 13139 20791
rect 13630 20788 13636 20800
rect 13127 20760 13636 20788
rect 13127 20757 13139 20760
rect 13081 20751 13139 20757
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14476 20788 14504 20816
rect 13872 20760 14504 20788
rect 13872 20748 13878 20760
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 16117 20791 16175 20797
rect 14884 20760 14929 20788
rect 14884 20748 14890 20760
rect 16117 20757 16129 20791
rect 16163 20788 16175 20791
rect 16666 20788 16672 20800
rect 16163 20760 16672 20788
rect 16163 20757 16175 20760
rect 16117 20751 16175 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 17678 20788 17684 20800
rect 17639 20760 17684 20788
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 19610 20748 19616 20800
rect 19668 20788 19674 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 19668 20760 19809 20788
rect 19668 20748 19674 20760
rect 19797 20757 19809 20760
rect 19843 20757 19855 20791
rect 20622 20788 20628 20800
rect 20583 20760 20628 20788
rect 19797 20751 19855 20757
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 1104 20698 21436 20720
rect 1104 20646 7727 20698
rect 7779 20646 7791 20698
rect 7843 20646 7855 20698
rect 7907 20646 7919 20698
rect 7971 20646 7983 20698
rect 8035 20646 14504 20698
rect 14556 20646 14568 20698
rect 14620 20646 14632 20698
rect 14684 20646 14696 20698
rect 14748 20646 14760 20698
rect 14812 20646 21436 20698
rect 1104 20624 21436 20646
rect 2314 20584 2320 20596
rect 2275 20556 2320 20584
rect 2314 20544 2320 20556
rect 2372 20544 2378 20596
rect 3697 20587 3755 20593
rect 3697 20553 3709 20587
rect 3743 20584 3755 20587
rect 4154 20584 4160 20596
rect 3743 20556 4160 20584
rect 3743 20553 3755 20556
rect 3697 20547 3755 20553
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 5408 20556 5580 20584
rect 5408 20544 5414 20556
rect 1489 20519 1547 20525
rect 1489 20485 1501 20519
rect 1535 20516 1547 20519
rect 3050 20516 3056 20528
rect 1535 20488 3056 20516
rect 1535 20485 1547 20488
rect 1489 20479 1547 20485
rect 3050 20476 3056 20488
rect 3108 20476 3114 20528
rect 3145 20519 3203 20525
rect 3145 20485 3157 20519
rect 3191 20516 3203 20519
rect 4246 20516 4252 20528
rect 3191 20488 4252 20516
rect 3191 20485 3203 20488
rect 3145 20479 3203 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 5437 20473 5495 20479
rect 5437 20470 5449 20473
rect 2222 20448 2228 20460
rect 2183 20420 2228 20448
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 2915 20420 3832 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 2682 20380 2688 20392
rect 1719 20352 2688 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 3145 20383 3203 20389
rect 3145 20380 3157 20383
rect 2884 20352 3157 20380
rect 2884 20324 2912 20352
rect 3145 20349 3157 20352
rect 3191 20349 3203 20383
rect 3804 20380 3832 20420
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 4617 20451 4675 20457
rect 3936 20420 3981 20448
rect 3936 20408 3942 20420
rect 4617 20417 4629 20451
rect 4663 20448 4675 20451
rect 4798 20448 4804 20460
rect 4663 20420 4804 20448
rect 4663 20417 4675 20420
rect 4617 20411 4675 20417
rect 4798 20408 4804 20420
rect 4856 20408 4862 20460
rect 5368 20442 5449 20470
rect 5368 20392 5396 20442
rect 5437 20439 5449 20442
rect 5483 20439 5495 20473
rect 5552 20457 5580 20556
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 6914 20584 6920 20596
rect 5960 20556 6920 20584
rect 5960 20544 5966 20556
rect 6914 20544 6920 20556
rect 6972 20584 6978 20596
rect 8110 20584 8116 20596
rect 6972 20556 8116 20584
rect 6972 20544 6978 20556
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 8662 20584 8668 20596
rect 8623 20556 8668 20584
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 10226 20584 10232 20596
rect 9824 20556 10232 20584
rect 9824 20544 9830 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 10870 20584 10876 20596
rect 10468 20556 10876 20584
rect 10468 20544 10474 20556
rect 10870 20544 10876 20556
rect 10928 20584 10934 20596
rect 10965 20587 11023 20593
rect 10965 20584 10977 20587
rect 10928 20556 10977 20584
rect 10928 20544 10934 20556
rect 10965 20553 10977 20556
rect 11011 20553 11023 20587
rect 10965 20547 11023 20553
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11572 20556 11621 20584
rect 11572 20544 11578 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 14553 20587 14611 20593
rect 11609 20547 11667 20553
rect 11716 20556 14504 20584
rect 5920 20516 5948 20544
rect 5721 20488 5948 20516
rect 5721 20457 5749 20488
rect 6270 20476 6276 20528
rect 6328 20516 6334 20528
rect 6549 20519 6607 20525
rect 6549 20516 6561 20519
rect 6328 20488 6561 20516
rect 6328 20476 6334 20488
rect 6549 20485 6561 20488
rect 6595 20516 6607 20519
rect 7282 20516 7288 20528
rect 6595 20488 7288 20516
rect 6595 20485 6607 20488
rect 6549 20479 6607 20485
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 7374 20476 7380 20528
rect 7432 20516 7438 20528
rect 8386 20516 8392 20528
rect 7432 20488 7880 20516
rect 7432 20476 7438 20488
rect 7852 20460 7880 20488
rect 7944 20488 8392 20516
rect 5437 20433 5495 20439
rect 5529 20451 5587 20457
rect 5529 20417 5541 20451
rect 5575 20417 5587 20451
rect 5529 20411 5587 20417
rect 5706 20451 5764 20457
rect 5706 20417 5718 20451
rect 5752 20417 5764 20451
rect 5706 20411 5764 20417
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 5868 20420 5913 20448
rect 5868 20408 5874 20420
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 6144 20420 6377 20448
rect 6144 20408 6150 20420
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6638 20448 6644 20460
rect 6599 20420 6644 20448
rect 6365 20411 6423 20417
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20417 6791 20451
rect 7650 20448 7656 20460
rect 7611 20420 7656 20448
rect 6733 20411 6791 20417
rect 4157 20383 4215 20389
rect 4157 20380 4169 20383
rect 3804 20352 4169 20380
rect 3145 20343 3203 20349
rect 4157 20349 4169 20352
rect 4203 20380 4215 20383
rect 4203 20352 4752 20380
rect 4203 20349 4215 20352
rect 4157 20343 4215 20349
rect 2866 20272 2872 20324
rect 2924 20272 2930 20324
rect 4724 20256 4752 20352
rect 5350 20340 5356 20392
rect 5408 20340 5414 20392
rect 6270 20340 6276 20392
rect 6328 20380 6334 20392
rect 6748 20380 6776 20411
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 7834 20448 7840 20460
rect 7747 20420 7840 20448
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 7944 20457 7972 20488
rect 8386 20476 8392 20488
rect 8444 20516 8450 20528
rect 8444 20488 8984 20516
rect 8444 20476 8450 20488
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20417 7987 20451
rect 8202 20448 8208 20460
rect 8163 20420 8208 20448
rect 7929 20411 7987 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8662 20448 8668 20460
rect 8623 20420 8668 20448
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 8754 20408 8760 20460
rect 8812 20448 8818 20460
rect 8956 20457 8984 20488
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 9732 20488 10180 20516
rect 9732 20476 9738 20488
rect 8849 20451 8907 20457
rect 8849 20448 8861 20451
rect 8812 20420 8861 20448
rect 8812 20408 8818 20420
rect 8849 20417 8861 20420
rect 8895 20417 8907 20451
rect 8849 20411 8907 20417
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9858 20448 9864 20460
rect 9819 20420 9864 20448
rect 9217 20411 9275 20417
rect 6328 20352 6776 20380
rect 6328 20340 6334 20352
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7742 20380 7748 20392
rect 7064 20352 7748 20380
rect 7064 20340 7070 20352
rect 7742 20340 7748 20352
rect 7800 20380 7806 20392
rect 9232 20380 9260 20411
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10152 20457 10180 20488
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20448 10195 20451
rect 10594 20448 10600 20460
rect 10183 20420 10600 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 7800 20352 9260 20380
rect 10060 20380 10088 20411
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 11606 20448 11612 20460
rect 11567 20420 11612 20448
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 10686 20380 10692 20392
rect 10060 20352 10692 20380
rect 7800 20340 7806 20352
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 11716 20380 11744 20556
rect 14093 20519 14151 20525
rect 11808 20488 13308 20516
rect 11808 20457 11836 20488
rect 13280 20460 13308 20488
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 14182 20516 14188 20528
rect 14139 20488 14188 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 14182 20476 14188 20488
rect 14240 20476 14246 20528
rect 14476 20516 14504 20556
rect 14553 20553 14565 20587
rect 14599 20584 14611 20587
rect 14826 20584 14832 20596
rect 14599 20556 14832 20584
rect 14599 20553 14611 20556
rect 14553 20547 14611 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15102 20544 15108 20596
rect 15160 20584 15166 20596
rect 15565 20587 15623 20593
rect 15565 20584 15577 20587
rect 15160 20556 15577 20584
rect 15160 20544 15166 20556
rect 15565 20553 15577 20556
rect 15611 20553 15623 20587
rect 15565 20547 15623 20553
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 16632 20556 16681 20584
rect 16632 20544 16638 20556
rect 16669 20553 16681 20556
rect 16715 20553 16727 20587
rect 17678 20584 17684 20596
rect 17639 20556 17684 20584
rect 16669 20547 16727 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 19242 20544 19248 20596
rect 19300 20584 19306 20596
rect 19797 20587 19855 20593
rect 19797 20584 19809 20587
rect 19300 20556 19809 20584
rect 19300 20544 19306 20556
rect 19797 20553 19809 20556
rect 19843 20553 19855 20587
rect 19797 20547 19855 20553
rect 16206 20516 16212 20528
rect 14476 20488 16212 20516
rect 16206 20476 16212 20488
rect 16264 20516 16270 20528
rect 16264 20488 16988 20516
rect 16264 20476 16270 20488
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 11900 20380 11928 20411
rect 11974 20408 11980 20460
rect 12032 20448 12038 20460
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 12032 20420 12173 20448
rect 12032 20408 12038 20420
rect 12161 20417 12173 20420
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12492 20420 12725 20448
rect 12492 20408 12498 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12894 20448 12900 20460
rect 12855 20420 12900 20448
rect 12713 20411 12771 20417
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 13262 20448 13268 20460
rect 13044 20420 13089 20448
rect 13223 20420 13268 20448
rect 13044 20408 13050 20420
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13906 20448 13912 20460
rect 13867 20420 13912 20448
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 14366 20408 14372 20460
rect 14424 20448 14430 20460
rect 14737 20451 14795 20457
rect 14737 20448 14749 20451
rect 14424 20420 14749 20448
rect 14424 20408 14430 20420
rect 14737 20417 14749 20420
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15102 20448 15108 20460
rect 14884 20420 14929 20448
rect 15063 20420 15108 20448
rect 14884 20408 14890 20420
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15344 20420 15761 20448
rect 15344 20408 15350 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 15654 20380 15660 20392
rect 11716 20352 11928 20380
rect 12360 20352 15660 20380
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 6178 20312 6184 20324
rect 5500 20284 6184 20312
rect 5500 20272 5506 20284
rect 6178 20272 6184 20284
rect 6236 20312 6242 20324
rect 6917 20315 6975 20321
rect 6917 20312 6929 20315
rect 6236 20284 6929 20312
rect 6236 20272 6242 20284
rect 6917 20281 6929 20284
rect 6963 20281 6975 20315
rect 6917 20275 6975 20281
rect 8021 20315 8079 20321
rect 8021 20281 8033 20315
rect 8067 20312 8079 20315
rect 8294 20312 8300 20324
rect 8067 20284 8300 20312
rect 8067 20281 8079 20284
rect 8021 20275 8079 20281
rect 8294 20272 8300 20284
rect 8352 20272 8358 20324
rect 9582 20272 9588 20324
rect 9640 20312 9646 20324
rect 9640 20284 10180 20312
rect 9640 20272 9646 20284
rect 2958 20244 2964 20256
rect 2919 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4065 20247 4123 20253
rect 4065 20244 4077 20247
rect 4028 20216 4077 20244
rect 4028 20204 4034 20216
rect 4065 20213 4077 20216
rect 4111 20213 4123 20247
rect 4706 20244 4712 20256
rect 4667 20216 4712 20244
rect 4065 20207 4123 20213
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 6822 20244 6828 20256
rect 5307 20216 6828 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 7650 20244 7656 20256
rect 7524 20216 7656 20244
rect 7524 20204 7530 20216
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8570 20244 8576 20256
rect 8159 20216 8576 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8570 20204 8576 20216
rect 8628 20244 8634 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8628 20216 9137 20244
rect 8628 20204 8634 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 9677 20247 9735 20253
rect 9677 20213 9689 20247
rect 9723 20244 9735 20247
rect 9950 20244 9956 20256
rect 9723 20216 9956 20244
rect 9723 20213 9735 20216
rect 9677 20207 9735 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10152 20244 10180 20284
rect 10226 20272 10232 20324
rect 10284 20312 10290 20324
rect 11808 20312 11836 20352
rect 10284 20284 11836 20312
rect 10284 20272 10290 20284
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 10152 20216 10609 20244
rect 10597 20213 10609 20216
rect 10643 20213 10655 20247
rect 10597 20207 10655 20213
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11020 20216 12081 20244
rect 11020 20204 11026 20216
rect 12069 20213 12081 20216
rect 12115 20244 12127 20247
rect 12360 20244 12388 20352
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 15764 20380 15792 20411
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16117 20451 16175 20457
rect 15896 20420 15941 20448
rect 15896 20408 15902 20420
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16390 20448 16396 20460
rect 16163 20420 16396 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 16960 20457 16988 20488
rect 17310 20476 17316 20528
rect 17368 20516 17374 20528
rect 17368 20488 17908 20516
rect 17368 20476 17374 20488
rect 17880 20457 17908 20488
rect 18506 20476 18512 20528
rect 18564 20516 18570 20528
rect 18601 20519 18659 20525
rect 18601 20516 18613 20519
rect 18564 20488 18613 20516
rect 18564 20476 18570 20488
rect 18601 20485 18613 20488
rect 18647 20485 18659 20519
rect 18601 20479 18659 20485
rect 20254 20476 20260 20528
rect 20312 20516 20318 20528
rect 20441 20519 20499 20525
rect 20441 20516 20453 20519
rect 20312 20488 20453 20516
rect 20312 20476 20318 20488
rect 20441 20485 20453 20488
rect 20487 20485 20499 20519
rect 20441 20479 20499 20485
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 17865 20451 17923 20457
rect 17267 20420 17632 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 16298 20380 16304 20392
rect 15764 20352 16304 20380
rect 16298 20340 16304 20352
rect 16356 20380 16362 20392
rect 16868 20380 16896 20411
rect 17604 20392 17632 20420
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 18782 20448 18788 20460
rect 18743 20420 18788 20448
rect 17865 20411 17923 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 19702 20448 19708 20460
rect 19663 20420 19708 20448
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 16356 20352 16896 20380
rect 16356 20340 16362 20352
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 18141 20383 18199 20389
rect 18141 20380 18153 20383
rect 17644 20352 18153 20380
rect 17644 20340 17650 20352
rect 18141 20349 18153 20352
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 13170 20312 13176 20324
rect 13131 20284 13176 20312
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 13354 20272 13360 20324
rect 13412 20312 13418 20324
rect 18049 20315 18107 20321
rect 18049 20312 18061 20315
rect 13412 20284 18061 20312
rect 13412 20272 13418 20284
rect 18049 20281 18061 20284
rect 18095 20281 18107 20315
rect 18049 20275 18107 20281
rect 15010 20244 15016 20256
rect 12115 20216 12388 20244
rect 14971 20216 15016 20244
rect 12115 20213 12127 20216
rect 12069 20207 12127 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 15746 20204 15752 20256
rect 15804 20244 15810 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15804 20216 16037 20244
rect 15804 20204 15810 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17129 20247 17187 20253
rect 17129 20244 17141 20247
rect 16632 20216 17141 20244
rect 16632 20204 16638 20216
rect 17129 20213 17141 20216
rect 17175 20213 17187 20247
rect 18966 20244 18972 20256
rect 18927 20216 18972 20244
rect 17129 20207 17187 20213
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 20128 20216 20545 20244
rect 20128 20204 20134 20216
rect 20533 20213 20545 20216
rect 20579 20213 20591 20247
rect 20533 20207 20591 20213
rect 1104 20154 21436 20176
rect 1104 20102 4338 20154
rect 4390 20102 4402 20154
rect 4454 20102 4466 20154
rect 4518 20102 4530 20154
rect 4582 20102 4594 20154
rect 4646 20102 11116 20154
rect 11168 20102 11180 20154
rect 11232 20102 11244 20154
rect 11296 20102 11308 20154
rect 11360 20102 11372 20154
rect 11424 20102 17893 20154
rect 17945 20102 17957 20154
rect 18009 20102 18021 20154
rect 18073 20102 18085 20154
rect 18137 20102 18149 20154
rect 18201 20102 21436 20154
rect 1104 20080 21436 20102
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 6454 20040 6460 20052
rect 4764 20012 6040 20040
rect 6415 20012 6460 20040
rect 4764 20000 4770 20012
rect 1670 19932 1676 19984
rect 1728 19932 1734 19984
rect 3789 19975 3847 19981
rect 3789 19941 3801 19975
rect 3835 19972 3847 19975
rect 5902 19972 5908 19984
rect 3835 19944 5908 19972
rect 3835 19941 3847 19944
rect 3789 19935 3847 19941
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 6012 19972 6040 20012
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 7009 20043 7067 20049
rect 7009 20009 7021 20043
rect 7055 20040 7067 20043
rect 8662 20040 8668 20052
rect 7055 20012 8668 20040
rect 7055 20009 7067 20012
rect 7009 20003 7067 20009
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 8846 20000 8852 20052
rect 8904 20040 8910 20052
rect 10873 20043 10931 20049
rect 10873 20040 10885 20043
rect 8904 20012 10885 20040
rect 8904 20000 8910 20012
rect 10873 20009 10885 20012
rect 10919 20009 10931 20043
rect 10873 20003 10931 20009
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13722 20040 13728 20052
rect 13403 20012 13728 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 15746 20040 15752 20052
rect 15707 20012 15752 20040
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16390 20040 16396 20052
rect 16080 20012 16396 20040
rect 16080 20000 16086 20012
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 17126 20040 17132 20052
rect 17087 20012 17132 20040
rect 17126 20000 17132 20012
rect 17184 20000 17190 20052
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18601 20043 18659 20049
rect 18601 20040 18613 20043
rect 18472 20012 18613 20040
rect 18472 20000 18478 20012
rect 18601 20009 18613 20012
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 8202 19972 8208 19984
rect 6012 19944 8208 19972
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 9493 19975 9551 19981
rect 9493 19941 9505 19975
rect 9539 19972 9551 19975
rect 11514 19972 11520 19984
rect 9539 19944 11520 19972
rect 9539 19941 9551 19944
rect 9493 19935 9551 19941
rect 11514 19932 11520 19944
rect 11572 19972 11578 19984
rect 11572 19944 11652 19972
rect 11572 19932 11578 19944
rect 1688 19904 1716 19932
rect 4338 19904 4344 19916
rect 1688 19876 2774 19904
rect 4299 19876 4344 19904
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2746 19836 2774 19876
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 7006 19904 7012 19916
rect 4580 19876 7012 19904
rect 4580 19864 4586 19876
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 7190 19864 7196 19916
rect 7248 19904 7254 19916
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 7248 19876 7389 19904
rect 7248 19864 7254 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19904 7527 19907
rect 7650 19904 7656 19916
rect 7515 19876 7656 19904
rect 7515 19873 7527 19876
rect 7469 19867 7527 19873
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8110 19864 8116 19916
rect 8168 19904 8174 19916
rect 8297 19907 8355 19913
rect 8297 19904 8309 19907
rect 8168 19876 8309 19904
rect 8168 19864 8174 19876
rect 8297 19873 8309 19876
rect 8343 19873 8355 19907
rect 9950 19904 9956 19916
rect 9911 19876 9956 19904
rect 8297 19867 8355 19873
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10042 19864 10048 19916
rect 10100 19904 10106 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 10100 19876 10149 19904
rect 10100 19864 10106 19876
rect 10137 19873 10149 19876
rect 10183 19904 10195 19907
rect 10778 19904 10784 19916
rect 10183 19876 10784 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 11624 19904 11652 19944
rect 11790 19932 11796 19984
rect 11848 19972 11854 19984
rect 14737 19975 14795 19981
rect 14737 19972 14749 19975
rect 11848 19944 14749 19972
rect 11848 19932 11854 19944
rect 14737 19941 14749 19944
rect 14783 19941 14795 19975
rect 14737 19935 14795 19941
rect 17957 19975 18015 19981
rect 17957 19941 17969 19975
rect 18003 19972 18015 19975
rect 18322 19972 18328 19984
rect 18003 19944 18328 19972
rect 18003 19941 18015 19944
rect 17957 19935 18015 19941
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 18230 19904 18236 19916
rect 11624 19876 12848 19904
rect 4706 19836 4712 19848
rect 2746 19808 4712 19836
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 5442 19836 5448 19848
rect 5403 19808 5448 19836
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5626 19836 5632 19848
rect 5587 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 7282 19836 7288 19848
rect 7243 19808 7288 19836
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19805 7619 19839
rect 7742 19836 7748 19848
rect 7703 19808 7748 19836
rect 7561 19799 7619 19805
rect 2866 19768 2872 19780
rect 2827 19740 2872 19768
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 3050 19768 3056 19780
rect 3011 19740 3056 19768
rect 3050 19728 3056 19740
rect 3108 19728 3114 19780
rect 6365 19771 6423 19777
rect 3252 19740 6316 19768
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 3252 19709 3280 19740
rect 3237 19703 3295 19709
rect 3237 19700 3249 19703
rect 3200 19672 3249 19700
rect 3200 19660 3206 19672
rect 3237 19669 3249 19672
rect 3283 19669 3295 19703
rect 3237 19663 3295 19669
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4157 19703 4215 19709
rect 4157 19700 4169 19703
rect 4120 19672 4169 19700
rect 4120 19660 4126 19672
rect 4157 19669 4169 19672
rect 4203 19669 4215 19703
rect 4157 19663 4215 19669
rect 4246 19660 4252 19712
rect 4304 19700 4310 19712
rect 4304 19672 4349 19700
rect 4304 19660 4310 19672
rect 5166 19660 5172 19712
rect 5224 19700 5230 19712
rect 5626 19700 5632 19712
rect 5224 19672 5632 19700
rect 5224 19660 5230 19672
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 5810 19700 5816 19712
rect 5771 19672 5816 19700
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 6288 19700 6316 19740
rect 6365 19737 6377 19771
rect 6411 19768 6423 19771
rect 6730 19768 6736 19780
rect 6411 19740 6736 19768
rect 6411 19737 6423 19740
rect 6365 19731 6423 19737
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 7576 19768 7604 19799
rect 7742 19796 7748 19808
rect 7800 19796 7806 19848
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 8202 19836 8208 19848
rect 7892 19808 8208 19836
rect 7892 19796 7898 19808
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 9306 19836 9312 19848
rect 8720 19808 9312 19836
rect 8720 19796 8726 19808
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 11425 19839 11483 19845
rect 11425 19836 11437 19839
rect 9640 19808 11437 19836
rect 9640 19796 9646 19808
rect 11425 19805 11437 19808
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12710 19836 12716 19848
rect 12575 19808 12716 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 12820 19845 12848 19876
rect 13096 19876 18236 19904
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 8110 19768 8116 19780
rect 7576 19740 8116 19768
rect 8110 19728 8116 19740
rect 8168 19768 8174 19780
rect 8478 19768 8484 19780
rect 8168 19740 8484 19768
rect 8168 19728 8174 19740
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 9030 19728 9036 19780
rect 9088 19768 9094 19780
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 9088 19740 10793 19768
rect 9088 19728 9094 19740
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 10781 19731 10839 19737
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 13096 19768 13124 19876
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 13262 19836 13268 19848
rect 13175 19808 13268 19836
rect 13262 19796 13268 19808
rect 13320 19836 13326 19848
rect 15470 19836 15476 19848
rect 13320 19808 15476 19836
rect 13320 19796 13326 19808
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 15838 19836 15844 19848
rect 15703 19808 15844 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 16298 19836 16304 19848
rect 16259 19808 16304 19836
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17276 19808 17785 19836
rect 17276 19796 17282 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 20438 19836 20444 19848
rect 20399 19808 20444 19836
rect 17773 19799 17831 19805
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 10928 19740 13124 19768
rect 10928 19728 10934 19740
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 14148 19740 14565 19768
rect 14148 19728 14154 19740
rect 14553 19737 14565 19740
rect 14599 19737 14611 19771
rect 15488 19768 15516 19796
rect 15930 19768 15936 19780
rect 15488 19740 15936 19768
rect 14553 19731 14611 19737
rect 15930 19728 15936 19740
rect 15988 19728 15994 19780
rect 17034 19768 17040 19780
rect 16995 19740 17040 19768
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 18509 19771 18567 19777
rect 18509 19737 18521 19771
rect 18555 19768 18567 19771
rect 18598 19768 18604 19780
rect 18555 19740 18604 19768
rect 18555 19737 18567 19740
rect 18509 19731 18567 19737
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 19794 19768 19800 19780
rect 19755 19740 19800 19768
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 9674 19700 9680 19712
rect 6288 19672 9680 19700
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 9858 19700 9864 19712
rect 9819 19672 9864 19700
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 11974 19700 11980 19712
rect 11563 19672 11980 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 12342 19700 12348 19712
rect 12303 19672 12348 19700
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 12710 19700 12716 19712
rect 12671 19672 12716 19700
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 16482 19700 16488 19712
rect 15712 19672 16488 19700
rect 15712 19660 15718 19672
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 19886 19700 19892 19712
rect 19847 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 1104 19610 21436 19632
rect 1104 19558 7727 19610
rect 7779 19558 7791 19610
rect 7843 19558 7855 19610
rect 7907 19558 7919 19610
rect 7971 19558 7983 19610
rect 8035 19558 14504 19610
rect 14556 19558 14568 19610
rect 14620 19558 14632 19610
rect 14684 19558 14696 19610
rect 14748 19558 14760 19610
rect 14812 19558 21436 19610
rect 1104 19536 21436 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 2961 19499 3019 19505
rect 2961 19465 2973 19499
rect 3007 19496 3019 19499
rect 3142 19496 3148 19508
rect 3007 19468 3148 19496
rect 3007 19465 3019 19468
rect 2961 19459 3019 19465
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 4062 19496 4068 19508
rect 4023 19468 4068 19496
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 5077 19499 5135 19505
rect 5077 19465 5089 19499
rect 5123 19496 5135 19499
rect 5718 19496 5724 19508
rect 5123 19468 5724 19496
rect 5123 19465 5135 19468
rect 5077 19459 5135 19465
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 8662 19496 8668 19508
rect 6472 19468 8668 19496
rect 3878 19388 3884 19440
rect 3936 19428 3942 19440
rect 5902 19428 5908 19440
rect 3936 19400 5580 19428
rect 3936 19388 3942 19400
rect 1486 19360 1492 19372
rect 1447 19332 1492 19360
rect 1486 19320 1492 19332
rect 1544 19320 1550 19372
rect 1670 19360 1676 19372
rect 1596 19332 1676 19360
rect 1210 19252 1216 19304
rect 1268 19292 1274 19304
rect 1596 19292 1624 19332
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 2130 19360 2136 19372
rect 2091 19332 2136 19360
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 2314 19360 2320 19372
rect 2275 19332 2320 19360
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 4264 19369 4292 19400
rect 3421 19363 3479 19369
rect 3421 19360 3433 19363
rect 2884 19332 3433 19360
rect 2884 19304 2912 19332
rect 3421 19329 3433 19332
rect 3467 19329 3479 19363
rect 3421 19323 3479 19329
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 4522 19360 4528 19372
rect 4483 19332 4528 19360
rect 4249 19323 4307 19329
rect 4522 19320 4528 19332
rect 4580 19320 4586 19372
rect 4982 19360 4988 19372
rect 4943 19332 4988 19360
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 1268 19264 1624 19292
rect 2501 19295 2559 19301
rect 1268 19252 1274 19264
rect 2501 19261 2513 19295
rect 2547 19292 2559 19295
rect 2866 19292 2872 19304
rect 2547 19264 2872 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3329 19295 3387 19301
rect 3329 19292 3341 19295
rect 3108 19264 3341 19292
rect 3108 19252 3114 19264
rect 3329 19261 3341 19264
rect 3375 19292 3387 19295
rect 3786 19292 3792 19304
rect 3375 19264 3792 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4540 19292 4568 19320
rect 4212 19264 4568 19292
rect 5552 19292 5580 19400
rect 5644 19400 5908 19428
rect 5644 19369 5672 19400
rect 5902 19388 5908 19400
rect 5960 19428 5966 19440
rect 6270 19428 6276 19440
rect 5960 19400 6276 19428
rect 5960 19388 5966 19400
rect 6270 19388 6276 19400
rect 6328 19388 6334 19440
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19329 5687 19363
rect 6472 19360 6500 19468
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 9033 19499 9091 19505
rect 9033 19465 9045 19499
rect 9079 19496 9091 19499
rect 9858 19496 9864 19508
rect 9079 19468 9864 19496
rect 9079 19465 9091 19468
rect 9033 19459 9091 19465
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 13078 19496 13084 19508
rect 13039 19468 13084 19496
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13780 19468 14136 19496
rect 13780 19456 13786 19468
rect 6733 19431 6791 19437
rect 6733 19397 6745 19431
rect 6779 19428 6791 19431
rect 7006 19428 7012 19440
rect 6779 19400 7012 19428
rect 6779 19397 6791 19400
rect 6733 19391 6791 19397
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 8389 19431 8447 19437
rect 8389 19428 8401 19431
rect 7300 19400 8401 19428
rect 7300 19372 7328 19400
rect 8389 19397 8401 19400
rect 8435 19397 8447 19431
rect 8389 19391 8447 19397
rect 8478 19388 8484 19440
rect 8536 19428 8542 19440
rect 8536 19400 9444 19428
rect 8536 19388 8542 19400
rect 6638 19360 6644 19372
rect 5629 19323 5687 19329
rect 5736 19332 6500 19360
rect 6599 19332 6644 19360
rect 5736 19292 5764 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 6822 19360 6828 19372
rect 6783 19332 6828 19360
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19360 7159 19363
rect 7282 19360 7288 19372
rect 7147 19332 7288 19360
rect 7147 19329 7159 19332
rect 7101 19323 7159 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7650 19360 7656 19372
rect 7611 19332 7656 19360
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8754 19360 8760 19372
rect 8343 19332 8760 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8754 19320 8760 19332
rect 8812 19360 8818 19372
rect 9122 19360 9128 19372
rect 8812 19332 9128 19360
rect 8812 19320 8818 19332
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9306 19360 9312 19372
rect 9263 19332 9312 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 9416 19369 9444 19400
rect 9508 19400 10548 19428
rect 9508 19369 9536 19400
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9766 19360 9772 19372
rect 9493 19323 9551 19329
rect 9600 19332 9772 19360
rect 5552 19264 5764 19292
rect 9416 19292 9444 19323
rect 9600 19292 9628 19332
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 9950 19360 9956 19372
rect 9911 19332 9956 19360
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 10134 19360 10140 19372
rect 10095 19332 10140 19360
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 10520 19369 10548 19400
rect 11698 19388 11704 19440
rect 11756 19428 11762 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 11756 19400 12173 19428
rect 11756 19388 11762 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 12253 19431 12311 19437
rect 12253 19397 12265 19431
rect 12299 19428 12311 19431
rect 12710 19428 12716 19440
rect 12299 19400 12716 19428
rect 12299 19397 12311 19400
rect 12253 19391 12311 19397
rect 10505 19363 10563 19369
rect 10284 19332 10329 19360
rect 10284 19320 10290 19332
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 10594 19360 10600 19372
rect 10551 19332 10600 19360
rect 10551 19329 10563 19332
rect 10505 19323 10563 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 11974 19360 11980 19372
rect 11935 19332 11980 19360
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12268 19360 12296 19391
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 12802 19388 12808 19440
rect 12860 19428 12866 19440
rect 13354 19428 13360 19440
rect 12860 19400 13360 19428
rect 12860 19388 12866 19400
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13998 19428 14004 19440
rect 13959 19400 14004 19428
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 12124 19332 12296 19360
rect 12345 19363 12403 19369
rect 12124 19320 12130 19332
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 13170 19360 13176 19372
rect 13035 19332 13176 19360
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 9416 19264 9628 19292
rect 10413 19295 10471 19301
rect 4212 19252 4218 19264
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 10962 19292 10968 19304
rect 10459 19264 10968 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11514 19252 11520 19304
rect 11572 19292 11578 19304
rect 12360 19292 12388 19323
rect 13170 19320 13176 19332
rect 13228 19360 13234 19372
rect 14108 19369 14136 19468
rect 15746 19456 15752 19508
rect 15804 19456 15810 19508
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 20625 19499 20683 19505
rect 20625 19496 20637 19499
rect 16356 19468 20637 19496
rect 16356 19456 16362 19468
rect 20625 19465 20637 19468
rect 20671 19465 20683 19499
rect 20625 19459 20683 19465
rect 15764 19428 15792 19456
rect 15764 19400 16160 19428
rect 14093 19363 14151 19369
rect 13228 19332 14044 19360
rect 13228 19320 13234 19332
rect 11572 19264 12388 19292
rect 11572 19252 11578 19264
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 13909 19295 13967 19301
rect 13909 19292 13921 19295
rect 13872 19264 13921 19292
rect 13872 19252 13878 19264
rect 13909 19261 13921 19264
rect 13955 19261 13967 19295
rect 14016 19292 14044 19332
rect 14093 19329 14105 19363
rect 14139 19329 14151 19363
rect 14093 19323 14151 19329
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14240 19332 14841 19360
rect 14240 19320 14246 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 15470 19360 15476 19372
rect 14829 19323 14887 19329
rect 14936 19332 15476 19360
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 14016 19264 14289 19292
rect 13909 19255 13967 19261
rect 14277 19261 14289 19264
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 14936 19292 14964 19332
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 14415 19264 14964 19292
rect 15764 19292 15792 19323
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16022 19360 16028 19372
rect 15896 19332 15941 19360
rect 15983 19332 16028 19360
rect 15896 19320 15902 19332
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16132 19369 16160 19400
rect 17494 19388 17500 19440
rect 17552 19428 17558 19440
rect 17552 19400 17908 19428
rect 17552 19388 17558 19400
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16666 19360 16672 19372
rect 16627 19332 16672 19360
rect 16117 19323 16175 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 17880 19369 17908 19400
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 19797 19431 19855 19437
rect 19797 19428 19809 19431
rect 19392 19400 19809 19428
rect 19392 19388 19398 19400
rect 19797 19397 19809 19400
rect 19843 19397 19855 19431
rect 19797 19391 19855 19397
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18564 19332 19073 19360
rect 18564 19320 18570 19332
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 19300 19332 20545 19360
rect 19300 19320 19306 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 18049 19295 18107 19301
rect 15764 19264 16804 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 3605 19227 3663 19233
rect 3605 19193 3617 19227
rect 3651 19224 3663 19227
rect 3878 19224 3884 19236
rect 3651 19196 3884 19224
rect 3651 19193 3663 19196
rect 3605 19187 3663 19193
rect 3878 19184 3884 19196
rect 3936 19184 3942 19236
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 6178 19224 6184 19236
rect 5592 19196 6184 19224
rect 5592 19184 5598 19196
rect 6178 19184 6184 19196
rect 6236 19184 6242 19236
rect 6365 19227 6423 19233
rect 6365 19193 6377 19227
rect 6411 19224 6423 19227
rect 12434 19224 12440 19236
rect 6411 19196 12440 19224
rect 6411 19193 6423 19196
rect 6365 19187 6423 19193
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 12529 19227 12587 19233
rect 12529 19193 12541 19227
rect 12575 19224 12587 19227
rect 12986 19224 12992 19236
rect 12575 19196 12992 19224
rect 12575 19193 12587 19196
rect 12529 19187 12587 19193
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 14093 19227 14151 19233
rect 14093 19193 14105 19227
rect 14139 19224 14151 19227
rect 15838 19224 15844 19236
rect 14139 19196 15844 19224
rect 14139 19193 14151 19196
rect 14093 19187 14151 19193
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 16776 19168 16804 19264
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18322 19292 18328 19304
rect 18095 19264 18328 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18322 19252 18328 19264
rect 18380 19292 18386 19304
rect 18966 19292 18972 19304
rect 18380 19264 18972 19292
rect 18380 19252 18386 19264
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19208 19264 19993 19292
rect 19208 19252 19214 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19224 19303 19227
rect 20806 19224 20812 19236
rect 19291 19196 20812 19224
rect 19291 19193 19303 19196
rect 19245 19187 19303 19193
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4120 19128 4445 19156
rect 4120 19116 4126 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 5721 19159 5779 19165
rect 5721 19125 5733 19159
rect 5767 19156 5779 19159
rect 6086 19156 6092 19168
rect 5767 19128 6092 19156
rect 5767 19125 5779 19128
rect 5721 19119 5779 19125
rect 6086 19116 6092 19128
rect 6144 19156 6150 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6144 19128 7021 19156
rect 6144 19116 6150 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 7098 19116 7104 19168
rect 7156 19156 7162 19168
rect 7745 19159 7803 19165
rect 7745 19156 7757 19159
rect 7156 19128 7757 19156
rect 7156 19116 7162 19128
rect 7745 19125 7757 19128
rect 7791 19125 7803 19159
rect 7745 19119 7803 19125
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 10284 19128 10333 19156
rect 10284 19116 10290 19128
rect 10321 19125 10333 19128
rect 10367 19125 10379 19159
rect 10321 19119 10379 19125
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 14182 19156 14188 19168
rect 12308 19128 14188 19156
rect 12308 19116 12314 19128
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14918 19156 14924 19168
rect 14879 19128 14924 19156
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 15565 19159 15623 19165
rect 15565 19125 15577 19159
rect 15611 19156 15623 19159
rect 15654 19156 15660 19168
rect 15611 19128 15660 19156
rect 15611 19125 15623 19128
rect 15565 19119 15623 19125
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 17957 19159 18015 19165
rect 17957 19125 17969 19159
rect 18003 19156 18015 19159
rect 18230 19156 18236 19168
rect 18003 19128 18236 19156
rect 18003 19125 18015 19128
rect 17957 19119 18015 19125
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 1104 19066 21436 19088
rect 1104 19014 4338 19066
rect 4390 19014 4402 19066
rect 4454 19014 4466 19066
rect 4518 19014 4530 19066
rect 4582 19014 4594 19066
rect 4646 19014 11116 19066
rect 11168 19014 11180 19066
rect 11232 19014 11244 19066
rect 11296 19014 11308 19066
rect 11360 19014 11372 19066
rect 11424 19014 17893 19066
rect 17945 19014 17957 19066
rect 18009 19014 18021 19066
rect 18073 19014 18085 19066
rect 18137 19014 18149 19066
rect 18201 19014 21436 19066
rect 1104 18992 21436 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 2222 18952 2228 18964
rect 1627 18924 2228 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 2958 18952 2964 18964
rect 2915 18924 2964 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4154 18952 4160 18964
rect 3927 18924 4160 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 5224 18924 5365 18952
rect 5224 18912 5230 18924
rect 5353 18921 5365 18924
rect 5399 18921 5411 18955
rect 5353 18915 5411 18921
rect 5813 18955 5871 18961
rect 5813 18921 5825 18955
rect 5859 18952 5871 18955
rect 6638 18952 6644 18964
rect 5859 18924 6644 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 8205 18955 8263 18961
rect 8205 18921 8217 18955
rect 8251 18952 8263 18955
rect 9030 18952 9036 18964
rect 8251 18924 9036 18952
rect 8251 18921 8263 18924
rect 8205 18915 8263 18921
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 11333 18955 11391 18961
rect 11333 18921 11345 18955
rect 11379 18952 11391 18955
rect 11974 18952 11980 18964
rect 11379 18924 11980 18952
rect 11379 18921 11391 18924
rect 11333 18915 11391 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 14182 18952 14188 18964
rect 14143 18924 14188 18952
rect 14182 18912 14188 18924
rect 14240 18952 14246 18964
rect 14918 18952 14924 18964
rect 14240 18924 14924 18952
rect 14240 18912 14246 18924
rect 14918 18912 14924 18924
rect 14976 18912 14982 18964
rect 16758 18952 16764 18964
rect 15580 18924 16764 18952
rect 1964 18856 6500 18884
rect 1964 18757 1992 18856
rect 2222 18816 2228 18828
rect 2183 18788 2228 18816
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18816 5595 18819
rect 5810 18816 5816 18828
rect 5583 18788 5816 18816
rect 5583 18785 5595 18788
rect 5537 18779 5595 18785
rect 5810 18776 5816 18788
rect 5868 18816 5874 18828
rect 6362 18816 6368 18828
rect 5868 18788 6368 18816
rect 5868 18776 5874 18788
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 6472 18816 6500 18856
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 9861 18887 9919 18893
rect 9861 18884 9873 18887
rect 6788 18856 9873 18884
rect 6788 18844 6794 18856
rect 9861 18853 9873 18856
rect 9907 18853 9919 18887
rect 9861 18847 9919 18853
rect 10318 18844 10324 18896
rect 10376 18884 10382 18896
rect 10376 18856 10548 18884
rect 10376 18844 10382 18856
rect 7282 18816 7288 18828
rect 6472 18788 7288 18816
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 10520 18825 10548 18856
rect 11514 18844 11520 18896
rect 11572 18884 11578 18896
rect 11885 18887 11943 18893
rect 11885 18884 11897 18887
rect 11572 18856 11897 18884
rect 11572 18844 11578 18856
rect 11885 18853 11897 18856
rect 11931 18853 11943 18887
rect 11885 18847 11943 18853
rect 12529 18887 12587 18893
rect 12529 18853 12541 18887
rect 12575 18884 12587 18887
rect 13354 18884 13360 18896
rect 12575 18856 13360 18884
rect 12575 18853 12587 18856
rect 12529 18847 12587 18853
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 10505 18819 10563 18825
rect 8404 18788 10364 18816
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2130 18708 2136 18760
rect 2188 18748 2194 18760
rect 2590 18748 2596 18760
rect 2188 18720 2596 18748
rect 2188 18708 2194 18720
rect 2590 18708 2596 18720
rect 2648 18748 2654 18760
rect 2777 18751 2835 18757
rect 2777 18748 2789 18751
rect 2648 18720 2789 18748
rect 2648 18708 2654 18720
rect 2777 18717 2789 18720
rect 2823 18717 2835 18751
rect 3786 18748 3792 18760
rect 3747 18720 3792 18748
rect 2777 18711 2835 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 3936 18720 4721 18748
rect 3936 18708 3942 18720
rect 4709 18717 4721 18720
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18717 5687 18751
rect 5629 18711 5687 18717
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18680 5411 18683
rect 5442 18680 5448 18692
rect 5399 18652 5448 18680
rect 5399 18649 5411 18652
rect 5353 18643 5411 18649
rect 5442 18640 5448 18652
rect 5500 18640 5506 18692
rect 5644 18680 5672 18711
rect 5902 18708 5908 18760
rect 5960 18748 5966 18760
rect 6457 18751 6515 18757
rect 6457 18748 6469 18751
rect 5960 18720 6469 18748
rect 5960 18708 5966 18720
rect 6457 18717 6469 18720
rect 6503 18748 6515 18751
rect 6730 18748 6736 18760
rect 6503 18720 6736 18748
rect 6503 18717 6515 18720
rect 6457 18711 6515 18717
rect 6730 18708 6736 18720
rect 6788 18708 6794 18760
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6845 18720 6929 18748
rect 5644 18652 5764 18680
rect 5736 18624 5764 18652
rect 5810 18640 5816 18692
rect 5868 18680 5874 18692
rect 6845 18680 6873 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7190 18708 7196 18760
rect 7248 18748 7254 18760
rect 8404 18757 8432 18788
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7248 18720 8401 18748
rect 7248 18708 7254 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 9030 18748 9036 18760
rect 8991 18720 9036 18748
rect 8389 18711 8447 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 10226 18748 10232 18760
rect 10187 18720 10232 18748
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10336 18748 10364 18788
rect 10505 18785 10517 18819
rect 10551 18816 10563 18819
rect 10778 18816 10784 18828
rect 10551 18788 10784 18816
rect 10551 18785 10563 18788
rect 10505 18779 10563 18785
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 12066 18816 12072 18828
rect 11992 18788 12072 18816
rect 10870 18748 10876 18760
rect 10336 18720 10876 18748
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11992 18757 12020 18788
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 13464 18788 14596 18816
rect 11458 18751 11516 18757
rect 11458 18748 11470 18751
rect 11440 18717 11470 18748
rect 11504 18748 11516 18751
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11504 18720 11989 18748
rect 11504 18717 11516 18720
rect 11440 18711 11516 18717
rect 11977 18717 11989 18720
rect 12023 18748 12035 18751
rect 12342 18748 12348 18760
rect 12023 18720 12348 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 5868 18652 6873 18680
rect 5868 18640 5874 18652
rect 10134 18640 10140 18692
rect 10192 18680 10198 18692
rect 11440 18680 11468 18711
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 12894 18748 12900 18760
rect 12855 18720 12900 18748
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 10192 18652 11468 18680
rect 10192 18640 10198 18652
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 13464 18680 13492 18788
rect 13998 18708 14004 18760
rect 14056 18748 14062 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 14056 18720 14105 18748
rect 14056 18708 14062 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14366 18748 14372 18760
rect 14327 18720 14372 18748
rect 14093 18711 14151 18717
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14568 18757 14596 18788
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 15470 18748 15476 18760
rect 15431 18720 15476 18748
rect 14553 18711 14611 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 15580 18757 15608 18924
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 17000 18924 17448 18952
rect 17000 18912 17006 18924
rect 16666 18884 16672 18896
rect 16579 18856 16672 18884
rect 15565 18751 15623 18757
rect 15565 18717 15577 18751
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 15712 18720 15757 18748
rect 15712 18708 15718 18720
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16482 18748 16488 18760
rect 15896 18720 15941 18748
rect 16443 18720 16488 18748
rect 15896 18708 15902 18720
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16592 18757 16620 18856
rect 16666 18844 16672 18856
rect 16724 18884 16730 18896
rect 17313 18887 17371 18893
rect 17313 18884 17325 18887
rect 16724 18856 17325 18884
rect 16724 18844 16730 18856
rect 17313 18853 17325 18856
rect 17359 18853 17371 18887
rect 17420 18884 17448 18924
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 17828 18924 18613 18952
rect 17828 18912 17834 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 18601 18915 18659 18921
rect 19613 18955 19671 18961
rect 19613 18921 19625 18955
rect 19659 18952 19671 18955
rect 19794 18952 19800 18964
rect 19659 18924 19800 18952
rect 19659 18921 19671 18924
rect 19613 18915 19671 18921
rect 19794 18912 19800 18924
rect 19852 18912 19858 18964
rect 17420 18856 19334 18884
rect 17313 18847 17371 18853
rect 17586 18776 17592 18828
rect 17644 18816 17650 18828
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 17644 18788 17877 18816
rect 17644 18776 17650 18788
rect 17865 18785 17877 18788
rect 17911 18785 17923 18819
rect 19306 18816 19334 18856
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 19306 18788 20269 18816
rect 17865 18779 17923 18785
rect 20257 18785 20269 18788
rect 20303 18816 20315 18819
rect 20622 18816 20628 18828
rect 20303 18788 20628 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16816 18720 16865 18748
rect 16816 18708 16822 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18748 17831 18751
rect 18230 18748 18236 18760
rect 17819 18720 18236 18748
rect 17819 18717 17831 18720
rect 17773 18711 17831 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18472 18720 18521 18748
rect 18472 18708 18478 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 18782 18748 18788 18760
rect 18555 18720 18788 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 12124 18652 13492 18680
rect 12124 18640 12130 18652
rect 15102 18640 15108 18692
rect 15160 18680 15166 18692
rect 16301 18683 16359 18689
rect 16301 18680 16313 18683
rect 15160 18652 16313 18680
rect 15160 18640 15166 18652
rect 16301 18649 16313 18652
rect 16347 18649 16359 18683
rect 16301 18643 16359 18649
rect 19794 18640 19800 18692
rect 19852 18680 19858 18692
rect 20073 18683 20131 18689
rect 20073 18680 20085 18683
rect 19852 18652 20085 18680
rect 19852 18640 19858 18652
rect 20073 18649 20085 18652
rect 20119 18649 20131 18683
rect 20073 18643 20131 18649
rect 2041 18615 2099 18621
rect 2041 18581 2053 18615
rect 2087 18612 2099 18615
rect 3418 18612 3424 18624
rect 2087 18584 3424 18612
rect 2087 18581 2099 18584
rect 2041 18575 2099 18581
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 4801 18615 4859 18621
rect 4801 18581 4813 18615
rect 4847 18612 4859 18615
rect 5626 18612 5632 18624
rect 4847 18584 5632 18612
rect 4847 18581 4859 18584
rect 4801 18575 4859 18581
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 5718 18572 5724 18624
rect 5776 18572 5782 18624
rect 6178 18572 6184 18624
rect 6236 18612 6242 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 6236 18584 6285 18612
rect 6236 18572 6242 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6273 18575 6331 18581
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 7101 18615 7159 18621
rect 7101 18612 7113 18615
rect 6972 18584 7113 18612
rect 6972 18572 6978 18584
rect 7101 18581 7113 18584
rect 7147 18581 7159 18615
rect 9122 18612 9128 18624
rect 9083 18584 9128 18612
rect 7101 18575 7159 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 10318 18612 10324 18624
rect 10279 18584 10324 18612
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 11514 18612 11520 18624
rect 11475 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12894 18612 12900 18624
rect 12308 18584 12900 18612
rect 12308 18572 12314 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 13044 18584 13089 18612
rect 13044 18572 13050 18584
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 14737 18615 14795 18621
rect 14737 18612 14749 18615
rect 14332 18584 14749 18612
rect 14332 18572 14338 18584
rect 14737 18581 14749 18584
rect 14783 18581 14795 18615
rect 14737 18575 14795 18581
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 15197 18615 15255 18621
rect 15197 18612 15209 18615
rect 14976 18584 15209 18612
rect 14976 18572 14982 18584
rect 15197 18581 15209 18584
rect 15243 18581 15255 18615
rect 17678 18612 17684 18624
rect 17639 18584 17684 18612
rect 15197 18575 15255 18581
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19981 18615 20039 18621
rect 19981 18612 19993 18615
rect 19392 18584 19993 18612
rect 19392 18572 19398 18584
rect 19981 18581 19993 18584
rect 20027 18581 20039 18615
rect 19981 18575 20039 18581
rect 1104 18522 21436 18544
rect 1104 18470 7727 18522
rect 7779 18470 7791 18522
rect 7843 18470 7855 18522
rect 7907 18470 7919 18522
rect 7971 18470 7983 18522
rect 8035 18470 14504 18522
rect 14556 18470 14568 18522
rect 14620 18470 14632 18522
rect 14684 18470 14696 18522
rect 14748 18470 14760 18522
rect 14812 18470 21436 18522
rect 1104 18448 21436 18470
rect 1670 18408 1676 18420
rect 1631 18380 1676 18408
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 2590 18408 2596 18420
rect 2551 18380 2596 18408
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 3418 18408 3424 18420
rect 3379 18380 3424 18408
rect 3418 18368 3424 18380
rect 3476 18368 3482 18420
rect 3513 18411 3571 18417
rect 3513 18377 3525 18411
rect 3559 18408 3571 18411
rect 5718 18408 5724 18420
rect 3559 18380 5724 18408
rect 3559 18377 3571 18380
rect 3513 18371 3571 18377
rect 2406 18340 2412 18352
rect 2367 18312 2412 18340
rect 2406 18300 2412 18312
rect 2464 18300 2470 18352
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 3237 18275 3295 18281
rect 2271 18244 3188 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3160 18204 3188 18244
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 3528 18272 3556 18371
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 6546 18408 6552 18420
rect 5859 18380 6552 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7006 18408 7012 18420
rect 6967 18380 7012 18408
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 10376 18380 11529 18408
rect 10376 18368 10382 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12986 18408 12992 18420
rect 12575 18380 12992 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 14366 18408 14372 18420
rect 14327 18380 14372 18408
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 15654 18368 15660 18420
rect 15712 18408 15718 18420
rect 16114 18408 16120 18420
rect 15712 18380 16120 18408
rect 15712 18368 15718 18380
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 17678 18408 17684 18420
rect 17175 18380 17684 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 19794 18408 19800 18420
rect 19755 18380 19800 18408
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20254 18408 20260 18420
rect 20027 18380 20260 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 5537 18343 5595 18349
rect 5537 18309 5549 18343
rect 5583 18340 5595 18343
rect 6733 18343 6791 18349
rect 6733 18340 6745 18343
rect 5583 18312 6745 18340
rect 5583 18309 5595 18312
rect 5537 18303 5595 18309
rect 6733 18309 6745 18312
rect 6779 18340 6791 18343
rect 7190 18340 7196 18352
rect 6779 18312 7196 18340
rect 6779 18309 6791 18312
rect 6733 18303 6791 18309
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 7929 18343 7987 18349
rect 7929 18340 7941 18343
rect 7340 18312 7941 18340
rect 7340 18300 7346 18312
rect 7929 18309 7941 18312
rect 7975 18309 7987 18343
rect 10594 18340 10600 18352
rect 10555 18312 10600 18340
rect 7929 18303 7987 18309
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 16206 18340 16212 18352
rect 16119 18312 16212 18340
rect 3283 18244 3556 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4065 18275 4123 18281
rect 4065 18272 4077 18275
rect 4028 18244 4077 18272
rect 4028 18232 4034 18244
rect 4065 18241 4077 18244
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 5074 18232 5080 18284
rect 5132 18272 5138 18284
rect 5261 18275 5319 18281
rect 5261 18272 5273 18275
rect 5132 18244 5273 18272
rect 5132 18232 5138 18244
rect 5261 18241 5273 18244
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 5445 18275 5503 18281
rect 5445 18272 5457 18275
rect 5408 18244 5457 18272
rect 5408 18232 5414 18244
rect 5445 18241 5457 18244
rect 5491 18241 5503 18275
rect 5626 18272 5632 18284
rect 5587 18244 5632 18272
rect 5445 18235 5503 18241
rect 3326 18204 3332 18216
rect 3160 18176 3332 18204
rect 3053 18167 3111 18173
rect 3068 18136 3096 18167
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18173 3663 18207
rect 5460 18204 5488 18235
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 6362 18272 6368 18284
rect 6323 18244 6368 18272
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6458 18275 6516 18281
rect 6458 18241 6470 18275
rect 6504 18241 6516 18275
rect 6638 18272 6644 18284
rect 6599 18244 6644 18272
rect 6458 18235 6516 18241
rect 6473 18204 6501 18235
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 6830 18275 6888 18281
rect 6830 18272 6842 18275
rect 6748 18244 6842 18272
rect 6546 18204 6552 18216
rect 5460 18176 6552 18204
rect 3605 18167 3663 18173
rect 3620 18136 3648 18167
rect 6546 18164 6552 18176
rect 6604 18164 6610 18216
rect 6748 18148 6776 18244
rect 6830 18241 6842 18244
rect 6876 18241 6888 18275
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 6830 18235 6888 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8294 18272 8300 18284
rect 8255 18244 8300 18272
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8628 18244 8677 18272
rect 8628 18232 8634 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18272 8907 18275
rect 9122 18272 9128 18284
rect 8895 18244 9128 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9272 18244 9689 18272
rect 9272 18232 9278 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 10376 18244 10517 18272
rect 10376 18232 10382 18244
rect 10505 18241 10517 18244
rect 10551 18272 10563 18275
rect 10686 18272 10692 18284
rect 10551 18244 10692 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 11974 18272 11980 18284
rect 11839 18244 11980 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12526 18272 12532 18284
rect 12115 18244 12532 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 8754 18204 8760 18216
rect 8435 18176 8760 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 9766 18204 9772 18216
rect 9727 18176 9772 18204
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 10042 18204 10048 18216
rect 9999 18176 10048 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 11716 18204 11744 18232
rect 11716 18176 12434 18204
rect 5534 18136 5540 18148
rect 3068 18108 5540 18136
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 6730 18136 6736 18148
rect 5684 18108 6736 18136
rect 5684 18096 5690 18108
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 11977 18139 12035 18145
rect 11977 18105 11989 18139
rect 12023 18136 12035 18139
rect 12066 18136 12072 18148
rect 12023 18108 12072 18136
rect 12023 18105 12035 18108
rect 11977 18099 12035 18105
rect 12066 18096 12072 18108
rect 12124 18096 12130 18148
rect 12406 18136 12434 18176
rect 12618 18136 12624 18148
rect 12406 18108 12624 18136
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 12728 18136 12756 18235
rect 12820 18204 12848 18235
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 12952 18244 13093 18272
rect 12952 18232 12958 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13170 18232 13176 18284
rect 13228 18272 13234 18284
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 13228 18244 13553 18272
rect 13228 18232 13234 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 13872 18244 14289 18272
rect 13872 18232 13878 18244
rect 14277 18241 14289 18244
rect 14323 18272 14335 18275
rect 15102 18272 15108 18284
rect 14323 18244 15108 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16022 18272 16028 18284
rect 15979 18244 16028 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16132 18281 16160 18312
rect 16206 18300 16212 18312
rect 16264 18340 16270 18352
rect 16264 18312 17632 18340
rect 16264 18300 16270 18312
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 17310 18272 17316 18284
rect 16632 18244 17316 18272
rect 16632 18232 16638 18244
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17604 18281 17632 18312
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18272 17647 18275
rect 17770 18272 17776 18284
rect 17635 18244 17776 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18272 18199 18275
rect 18782 18272 18788 18284
rect 18187 18244 18788 18272
rect 18187 18241 18199 18244
rect 18141 18235 18199 18241
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 19058 18272 19064 18284
rect 19019 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 19978 18272 19984 18284
rect 19939 18244 19984 18272
rect 19978 18232 19984 18244
rect 20036 18272 20042 18284
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 20036 18244 20453 18272
rect 20036 18232 20042 18244
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 13633 18207 13691 18213
rect 13633 18204 13645 18207
rect 12820 18176 13645 18204
rect 13633 18173 13645 18176
rect 13679 18173 13691 18207
rect 13633 18167 13691 18173
rect 15470 18164 15476 18216
rect 15528 18204 15534 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15528 18176 15669 18204
rect 15528 18164 15534 18176
rect 15657 18173 15669 18176
rect 15703 18204 15715 18207
rect 15746 18204 15752 18216
rect 15703 18176 15752 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 15746 18164 15752 18176
rect 15804 18204 15810 18216
rect 16758 18204 16764 18216
rect 15804 18176 16764 18204
rect 15804 18164 15810 18176
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 14182 18136 14188 18148
rect 12728 18108 14188 18136
rect 14182 18096 14188 18108
rect 14240 18096 14246 18148
rect 18690 18136 18696 18148
rect 14936 18108 18696 18136
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18068 4215 18071
rect 4246 18068 4252 18080
rect 4203 18040 4252 18068
rect 4203 18037 4215 18040
rect 4157 18031 4215 18037
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 7064 18040 9321 18068
rect 7064 18028 7070 18040
rect 9309 18037 9321 18040
rect 9355 18037 9367 18071
rect 9309 18031 9367 18037
rect 12989 18071 13047 18077
rect 12989 18037 13001 18071
rect 13035 18068 13047 18071
rect 13078 18068 13084 18080
rect 13035 18040 13084 18068
rect 13035 18037 13047 18040
rect 12989 18031 13047 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 14936 18068 14964 18108
rect 18690 18096 18696 18108
rect 18748 18096 18754 18148
rect 15378 18068 15384 18080
rect 13320 18040 14964 18068
rect 15339 18040 15384 18068
rect 13320 18028 13326 18040
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 15712 18040 15761 18068
rect 15712 18028 15718 18040
rect 15749 18037 15761 18040
rect 15795 18037 15807 18071
rect 15749 18031 15807 18037
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 15896 18040 15941 18068
rect 15896 18028 15902 18040
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16390 18068 16396 18080
rect 16080 18040 16396 18068
rect 16080 18028 16086 18040
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 17497 18071 17555 18077
rect 17497 18068 17509 18071
rect 17092 18040 17509 18068
rect 17092 18028 17098 18040
rect 17497 18037 17509 18040
rect 17543 18037 17555 18071
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 17497 18031 17555 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19245 18071 19303 18077
rect 19245 18068 19257 18071
rect 19024 18040 19257 18068
rect 19024 18028 19030 18040
rect 19245 18037 19257 18040
rect 19291 18037 19303 18071
rect 19245 18031 19303 18037
rect 20254 18028 20260 18080
rect 20312 18068 20318 18080
rect 20349 18071 20407 18077
rect 20349 18068 20361 18071
rect 20312 18040 20361 18068
rect 20312 18028 20318 18040
rect 20349 18037 20361 18040
rect 20395 18037 20407 18071
rect 20349 18031 20407 18037
rect 1104 17978 21436 18000
rect 1104 17926 4338 17978
rect 4390 17926 4402 17978
rect 4454 17926 4466 17978
rect 4518 17926 4530 17978
rect 4582 17926 4594 17978
rect 4646 17926 11116 17978
rect 11168 17926 11180 17978
rect 11232 17926 11244 17978
rect 11296 17926 11308 17978
rect 11360 17926 11372 17978
rect 11424 17926 17893 17978
rect 17945 17926 17957 17978
rect 18009 17926 18021 17978
rect 18073 17926 18085 17978
rect 18137 17926 18149 17978
rect 18201 17926 21436 17978
rect 1104 17904 21436 17926
rect 5445 17867 5503 17873
rect 5445 17833 5457 17867
rect 5491 17864 5503 17867
rect 5718 17864 5724 17876
rect 5491 17836 5724 17864
rect 5491 17833 5503 17836
rect 5445 17827 5503 17833
rect 5718 17824 5724 17836
rect 5776 17864 5782 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5776 17836 6469 17864
rect 5776 17824 5782 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 6546 17824 6552 17876
rect 6604 17864 6610 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 6604 17836 7389 17864
rect 6604 17824 6610 17836
rect 7377 17833 7389 17836
rect 7423 17833 7435 17867
rect 7377 17827 7435 17833
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 9214 17864 9220 17876
rect 7975 17836 9220 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 10686 17864 10692 17876
rect 9548 17836 10692 17864
rect 9548 17824 9554 17836
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 12066 17864 12072 17876
rect 12027 17836 12072 17864
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12676 17836 12725 17864
rect 12676 17824 12682 17836
rect 12713 17833 12725 17836
rect 12759 17833 12771 17867
rect 12713 17827 12771 17833
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 13722 17864 13728 17876
rect 13403 17836 13728 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 14332 17836 14473 17864
rect 14332 17824 14338 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 15105 17867 15163 17873
rect 15105 17864 15117 17867
rect 14884 17836 15117 17864
rect 14884 17824 14890 17836
rect 15105 17833 15117 17836
rect 15151 17833 15163 17867
rect 15105 17827 15163 17833
rect 15562 17824 15568 17876
rect 15620 17864 15626 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 15620 17836 15669 17864
rect 15620 17824 15626 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 15657 17827 15715 17833
rect 16022 17824 16028 17876
rect 16080 17864 16086 17876
rect 16298 17864 16304 17876
rect 16080 17836 16304 17864
rect 16080 17824 16086 17836
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 16758 17864 16764 17876
rect 16719 17836 16764 17864
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 18509 17867 18567 17873
rect 18509 17833 18521 17867
rect 18555 17864 18567 17867
rect 19334 17864 19340 17876
rect 18555 17836 19340 17864
rect 18555 17833 18567 17836
rect 18509 17827 18567 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 5258 17796 5264 17808
rect 4356 17768 5264 17796
rect 2406 17688 2412 17740
rect 2464 17728 2470 17740
rect 3970 17728 3976 17740
rect 2464 17700 3976 17728
rect 2464 17688 2470 17700
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 3068 17660 3096 17700
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4356 17737 4384 17768
rect 5258 17756 5264 17768
rect 5316 17756 5322 17808
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 8941 17799 8999 17805
rect 8941 17796 8953 17799
rect 7892 17768 8953 17796
rect 7892 17756 7898 17768
rect 8941 17765 8953 17768
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 9030 17756 9036 17808
rect 9088 17796 9094 17808
rect 9950 17796 9956 17808
rect 9088 17768 9444 17796
rect 9911 17768 9956 17796
rect 9088 17756 9094 17768
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 4212 17700 4353 17728
rect 4212 17688 4218 17700
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 8389 17731 8447 17737
rect 4341 17691 4399 17697
rect 5276 17700 6592 17728
rect 3145 17663 3203 17669
rect 3145 17660 3157 17663
rect 3068 17632 3157 17660
rect 3145 17629 3157 17632
rect 3191 17629 3203 17663
rect 3145 17623 3203 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3326 17660 3332 17672
rect 3283 17632 3332 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 5276 17669 5304 17700
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17629 5319 17663
rect 5534 17660 5540 17672
rect 5447 17632 5540 17660
rect 5261 17623 5319 17629
rect 5534 17620 5540 17632
rect 5592 17660 5598 17672
rect 5810 17660 5816 17672
rect 5592 17632 5816 17660
rect 5592 17620 5598 17632
rect 5810 17620 5816 17632
rect 5868 17620 5874 17672
rect 6178 17660 6184 17672
rect 6139 17632 6184 17660
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 6564 17669 6592 17700
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 8662 17728 8668 17740
rect 8435 17700 8668 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 8662 17688 8668 17700
rect 8720 17728 8726 17740
rect 9122 17728 9128 17740
rect 8720 17700 9128 17728
rect 8720 17688 8726 17700
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 9416 17737 9444 17768
rect 9950 17756 9956 17768
rect 10008 17756 10014 17808
rect 11517 17799 11575 17805
rect 10152 17768 10364 17796
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 10152 17728 10180 17768
rect 9447 17700 10180 17728
rect 10229 17731 10287 17737
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10336 17728 10364 17768
rect 11517 17765 11529 17799
rect 11563 17796 11575 17799
rect 18414 17796 18420 17808
rect 11563 17768 18420 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 18414 17756 18420 17768
rect 18472 17756 18478 17808
rect 18601 17799 18659 17805
rect 18601 17765 18613 17799
rect 18647 17796 18659 17799
rect 19518 17796 19524 17808
rect 18647 17768 19524 17796
rect 18647 17765 18659 17768
rect 18601 17759 18659 17765
rect 19518 17756 19524 17768
rect 19576 17756 19582 17808
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20438 17796 20444 17808
rect 20027 17768 20444 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 20438 17756 20444 17768
rect 20496 17796 20502 17808
rect 20533 17799 20591 17805
rect 20533 17796 20545 17799
rect 20496 17768 20545 17796
rect 20496 17756 20502 17768
rect 20533 17765 20545 17768
rect 20579 17765 20591 17799
rect 20533 17759 20591 17765
rect 10336 17700 12388 17728
rect 10229 17691 10287 17697
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17629 6423 17663
rect 6365 17623 6423 17629
rect 6549 17663 6607 17669
rect 6549 17629 6561 17663
rect 6595 17660 6607 17663
rect 6638 17660 6644 17672
rect 6595 17632 6644 17660
rect 6595 17629 6607 17632
rect 6549 17623 6607 17629
rect 1854 17592 1860 17604
rect 1815 17564 1860 17592
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 2777 17595 2835 17601
rect 2777 17561 2789 17595
rect 2823 17592 2835 17595
rect 4249 17595 4307 17601
rect 4249 17592 4261 17595
rect 2823 17564 4261 17592
rect 2823 17561 2835 17564
rect 2777 17555 2835 17561
rect 4249 17561 4261 17564
rect 4295 17561 4307 17595
rect 4249 17555 4307 17561
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 3789 17527 3847 17533
rect 3789 17493 3801 17527
rect 3835 17524 3847 17527
rect 3878 17524 3884 17536
rect 3835 17496 3884 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 4154 17524 4160 17536
rect 4115 17496 4160 17524
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 5074 17524 5080 17536
rect 5035 17496 5080 17524
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 6380 17524 6408 17623
rect 6638 17620 6644 17632
rect 6696 17620 6702 17672
rect 6730 17620 6736 17672
rect 6788 17660 6794 17672
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 6788 17632 7021 17660
rect 6788 17620 6794 17632
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7190 17660 7196 17672
rect 7151 17632 7196 17660
rect 7009 17623 7067 17629
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 7616 17632 8125 17660
rect 7616 17620 7622 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8478 17660 8484 17672
rect 8343 17632 8484 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8754 17620 8760 17672
rect 8812 17660 8818 17672
rect 9030 17660 9036 17672
rect 8812 17632 9036 17660
rect 8812 17620 8818 17632
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9490 17660 9496 17672
rect 9451 17632 9496 17660
rect 9217 17623 9275 17629
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 8772 17592 8800 17620
rect 9232 17592 9260 17623
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10134 17660 10140 17672
rect 10091 17632 10140 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10244 17604 10272 17691
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10376 17632 10425 17660
rect 10376 17620 10382 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10686 17660 10692 17672
rect 10551 17632 10692 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 11330 17660 11336 17672
rect 11291 17632 11336 17660
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 10226 17592 10232 17604
rect 6880 17564 8800 17592
rect 8956 17564 10232 17592
rect 6880 17552 6886 17564
rect 6840 17524 6868 17552
rect 6380 17496 6868 17524
rect 8478 17484 8484 17536
rect 8536 17524 8542 17536
rect 8956 17524 8984 17564
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 10594 17552 10600 17604
rect 10652 17592 10658 17604
rect 12360 17592 12388 17700
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 12710 17728 12716 17740
rect 12492 17700 12716 17728
rect 12492 17688 12498 17700
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 13998 17688 14004 17740
rect 14056 17728 14062 17740
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 14056 17700 14105 17728
rect 14056 17688 14062 17700
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14918 17728 14924 17740
rect 14093 17691 14151 17697
rect 14292 17700 14924 17728
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12584 17632 12633 17660
rect 12584 17620 12590 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 13630 17660 13636 17672
rect 13587 17632 13636 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 12636 17592 12664 17623
rect 13630 17620 13636 17632
rect 13688 17620 13694 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14292 17669 14320 17700
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 16114 17728 16120 17740
rect 16027 17700 16120 17728
rect 16114 17688 16120 17700
rect 16172 17728 16178 17740
rect 16574 17728 16580 17740
rect 16172 17700 16580 17728
rect 16172 17688 16178 17700
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 17184 17700 19334 17728
rect 17184 17688 17190 17700
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13872 17632 14289 17660
rect 13872 17620 13878 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 15010 17660 15016 17672
rect 14971 17632 15016 17660
rect 14553 17623 14611 17629
rect 14568 17592 14596 17623
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15378 17620 15384 17672
rect 15436 17660 15442 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15436 17632 15669 17660
rect 15436 17620 15442 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16022 17660 16028 17672
rect 15979 17632 16028 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 10652 17564 12204 17592
rect 12360 17564 12572 17592
rect 12636 17564 14596 17592
rect 10652 17552 10658 17564
rect 8536 17496 8984 17524
rect 9125 17527 9183 17533
rect 8536 17484 8542 17496
rect 9125 17493 9137 17527
rect 9171 17524 9183 17527
rect 9306 17524 9312 17536
rect 9171 17496 9312 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9306 17484 9312 17496
rect 9364 17524 9370 17536
rect 10137 17527 10195 17533
rect 10137 17524 10149 17527
rect 9364 17496 10149 17524
rect 9364 17484 9370 17496
rect 10137 17493 10149 17496
rect 10183 17493 10195 17527
rect 12176 17524 12204 17564
rect 12434 17524 12440 17536
rect 12176 17496 12440 17524
rect 10137 17487 10195 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12544 17524 12572 17564
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 15856 17592 15884 17623
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 16206 17660 16212 17672
rect 16167 17632 16212 17660
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16942 17660 16948 17672
rect 16715 17632 16948 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16482 17592 16488 17604
rect 15620 17564 16488 17592
rect 15620 17552 15626 17564
rect 16482 17552 16488 17564
rect 16540 17592 16546 17604
rect 16684 17592 16712 17623
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17660 17371 17663
rect 18138 17660 18144 17672
rect 17359 17632 18000 17660
rect 18099 17632 18144 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 16540 17564 16712 17592
rect 17497 17595 17555 17601
rect 16540 17552 16546 17564
rect 17497 17561 17509 17595
rect 17543 17592 17555 17595
rect 17972 17592 18000 17632
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 18340 17669 18368 17700
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18690 17660 18696 17672
rect 18472 17632 18517 17660
rect 18651 17632 18696 17660
rect 18472 17620 18478 17632
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19306 17660 19334 17700
rect 19904 17700 20760 17728
rect 19554 17663 19612 17669
rect 19554 17660 19566 17663
rect 19306 17632 19566 17660
rect 19554 17629 19566 17632
rect 19600 17660 19612 17663
rect 19904 17660 19932 17700
rect 19600 17632 19932 17660
rect 19600 17629 19612 17632
rect 19554 17623 19612 17629
rect 19978 17620 19984 17672
rect 20036 17660 20042 17672
rect 20073 17663 20131 17669
rect 20073 17660 20085 17663
rect 20036 17632 20085 17660
rect 20036 17620 20042 17632
rect 20073 17629 20085 17632
rect 20119 17629 20131 17663
rect 20530 17660 20536 17672
rect 20073 17623 20131 17629
rect 20177 17632 20536 17660
rect 18782 17592 18788 17604
rect 17543 17564 17908 17592
rect 17972 17564 18788 17592
rect 17543 17561 17555 17564
rect 17497 17555 17555 17561
rect 17512 17524 17540 17555
rect 12544 17496 17540 17524
rect 17681 17527 17739 17533
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 17770 17524 17776 17536
rect 17727 17496 17776 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 17880 17524 17908 17564
rect 18782 17552 18788 17564
rect 18840 17552 18846 17604
rect 19334 17592 19340 17604
rect 19306 17552 19340 17592
rect 19392 17552 19398 17604
rect 20177 17592 20205 17632
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 20732 17669 20760 17700
rect 20717 17663 20775 17669
rect 20717 17660 20729 17663
rect 20680 17632 20729 17660
rect 20680 17620 20686 17632
rect 20717 17629 20729 17632
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 19628 17564 20205 17592
rect 19306 17524 19334 17552
rect 19628 17536 19656 17564
rect 19426 17524 19432 17536
rect 17880 17496 19334 17524
rect 19387 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19610 17524 19616 17536
rect 19571 17496 19616 17524
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 1104 17434 21436 17456
rect 1104 17382 7727 17434
rect 7779 17382 7791 17434
rect 7843 17382 7855 17434
rect 7907 17382 7919 17434
rect 7971 17382 7983 17434
rect 8035 17382 14504 17434
rect 14556 17382 14568 17434
rect 14620 17382 14632 17434
rect 14684 17382 14696 17434
rect 14748 17382 14760 17434
rect 14812 17382 21436 17434
rect 1104 17360 21436 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 1765 17323 1823 17329
rect 1765 17320 1777 17323
rect 1636 17292 1777 17320
rect 1636 17280 1642 17292
rect 1765 17289 1777 17292
rect 1811 17289 1823 17323
rect 2498 17320 2504 17332
rect 2459 17292 2504 17320
rect 1765 17283 1823 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 3605 17323 3663 17329
rect 3605 17289 3617 17323
rect 3651 17320 3663 17323
rect 4154 17320 4160 17332
rect 3651 17292 4160 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5132 17292 5273 17320
rect 5132 17280 5138 17292
rect 5261 17289 5273 17292
rect 5307 17320 5319 17323
rect 6546 17320 6552 17332
rect 5307 17292 5672 17320
rect 6507 17292 6552 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 5534 17252 5540 17264
rect 2700 17224 5540 17252
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17184 2007 17187
rect 2038 17184 2044 17196
rect 1995 17156 2044 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 2038 17144 2044 17156
rect 2096 17184 2102 17196
rect 2700 17193 2728 17224
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 2096 17156 2697 17184
rect 2096 17144 2102 17156
rect 2685 17153 2697 17156
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 3694 17144 3700 17196
rect 3752 17184 3758 17196
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 3752 17156 3801 17184
rect 3752 17144 3758 17156
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4246 17184 4252 17196
rect 4111 17156 4252 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 5644 17193 5672 17292
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7006 17280 7012 17332
rect 7064 17280 7070 17332
rect 8941 17323 8999 17329
rect 7116 17292 8892 17320
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 7024 17252 7052 17280
rect 6236 17224 7052 17252
rect 6236 17212 6242 17224
rect 6380 17193 6408 17224
rect 5258 17187 5316 17193
rect 5258 17153 5270 17187
rect 5304 17153 5316 17187
rect 5258 17147 5316 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6822 17184 6828 17196
rect 6595 17156 6828 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 3973 17051 4031 17057
rect 3973 17017 3985 17051
rect 4019 17048 4031 17051
rect 4062 17048 4068 17060
rect 4019 17020 4068 17048
rect 4019 17017 4031 17020
rect 3973 17011 4031 17017
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 4264 17048 4292 17144
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5276 17116 5304 17147
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 7006 17184 7012 17196
rect 6967 17156 7012 17184
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 5224 17088 5733 17116
rect 5224 17076 5230 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 7116 17116 7144 17292
rect 8294 17252 8300 17264
rect 7300 17224 8300 17252
rect 7300 17193 7328 17224
rect 8294 17212 8300 17224
rect 8352 17252 8358 17264
rect 8754 17252 8760 17264
rect 8352 17224 8760 17252
rect 8352 17212 8358 17224
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 8864 17252 8892 17292
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 9766 17320 9772 17332
rect 8987 17292 9772 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 13262 17320 13268 17332
rect 11388 17292 13268 17320
rect 11388 17280 11394 17292
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 13909 17323 13967 17329
rect 13909 17320 13921 17323
rect 13504 17292 13921 17320
rect 13504 17280 13510 17292
rect 13909 17289 13921 17292
rect 13955 17289 13967 17323
rect 13909 17283 13967 17289
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14274 17320 14280 17332
rect 14056 17292 14280 17320
rect 14056 17280 14062 17292
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 14424 17292 14469 17320
rect 14424 17280 14430 17292
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 20070 17320 20076 17332
rect 14884 17292 20076 17320
rect 14884 17280 14890 17292
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 20254 17320 20260 17332
rect 20215 17292 20260 17320
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 20622 17320 20628 17332
rect 20583 17292 20628 17320
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 11974 17252 11980 17264
rect 8864 17224 9076 17252
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 8662 17184 8668 17196
rect 8623 17156 8668 17184
rect 7561 17147 7619 17153
rect 5868 17088 7144 17116
rect 7208 17116 7236 17147
rect 7374 17116 7380 17128
rect 7208 17088 7380 17116
rect 5868 17076 5874 17088
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 7576 17116 7604 17147
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 7524 17088 7604 17116
rect 7524 17076 7530 17088
rect 7576 17048 7604 17088
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 8904 17088 8953 17116
rect 8904 17076 8910 17088
rect 8941 17085 8953 17088
rect 8987 17085 8999 17119
rect 9048 17116 9076 17224
rect 9416 17224 11980 17252
rect 9416 17193 9444 17224
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 19426 17252 19432 17264
rect 12084 17224 19432 17252
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17184 10103 17187
rect 10594 17184 10600 17196
rect 10091 17156 10600 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10744 17156 10789 17184
rect 10744 17144 10750 17156
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11698 17184 11704 17196
rect 10928 17156 11704 17184
rect 10928 17144 10934 17156
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12084 17184 12112 17224
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 11993 17156 12112 17184
rect 12161 17187 12219 17193
rect 11993 17116 12021 17156
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17184 12955 17187
rect 14182 17184 14188 17196
rect 12943 17156 14188 17184
rect 12943 17153 12955 17156
rect 12897 17147 12955 17153
rect 9048 17088 12021 17116
rect 8941 17079 8999 17085
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12176 17116 12204 17147
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17182 14335 17187
rect 15286 17184 15292 17196
rect 14476 17182 15292 17184
rect 14323 17156 15292 17182
rect 14323 17154 14504 17156
rect 14323 17153 14335 17154
rect 14277 17147 14335 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15562 17184 15568 17196
rect 15436 17156 15481 17184
rect 15523 17156 15568 17184
rect 15436 17144 15442 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17184 15715 17187
rect 15930 17184 15936 17196
rect 15703 17156 15936 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17313 17190 17371 17193
rect 17052 17187 17371 17190
rect 17052 17184 17325 17187
rect 16632 17162 17325 17184
rect 16632 17156 17080 17162
rect 16632 17144 16638 17156
rect 17313 17153 17325 17162
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17405 17187 17463 17193
rect 17405 17153 17417 17187
rect 17451 17184 17463 17187
rect 17494 17184 17500 17196
rect 17451 17156 17500 17184
rect 17451 17153 17463 17156
rect 17405 17147 17463 17153
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 17678 17184 17684 17196
rect 17639 17156 17684 17184
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17184 18475 17187
rect 18506 17184 18512 17196
rect 18463 17156 18512 17184
rect 18463 17153 18475 17156
rect 18417 17147 18475 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17184 18659 17187
rect 18874 17184 18880 17196
rect 18647 17156 18880 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 19702 17184 19708 17196
rect 19567 17156 19708 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 20438 17184 20444 17196
rect 20399 17156 20444 17184
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20588 17156 20729 17184
rect 20588 17144 20594 17156
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 12124 17088 12204 17116
rect 12124 17076 12130 17088
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 13228 17088 14473 17116
rect 13228 17076 13234 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 17126 17116 17132 17128
rect 16724 17088 17132 17116
rect 16724 17076 16730 17088
rect 17126 17076 17132 17088
rect 17184 17116 17190 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17184 17088 17233 17116
rect 17184 17076 17190 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 18138 17116 18144 17128
rect 17221 17079 17279 17085
rect 17420 17088 18144 17116
rect 4264 17020 7604 17048
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 13998 17048 14004 17060
rect 8803 17020 14004 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 17420 17057 17448 17088
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 18748 17088 19809 17116
rect 18748 17076 18754 17088
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 19797 17079 19855 17085
rect 17405 17051 17463 17057
rect 17405 17017 17417 17051
rect 17451 17017 17463 17051
rect 18782 17048 18788 17060
rect 18743 17020 18788 17048
rect 17405 17011 17463 17017
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 5077 16983 5135 16989
rect 5077 16949 5089 16983
rect 5123 16980 5135 16983
rect 6362 16980 6368 16992
rect 5123 16952 6368 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 7009 16983 7067 16989
rect 7009 16949 7021 16983
rect 7055 16980 7067 16983
rect 7098 16980 7104 16992
rect 7055 16952 7104 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7469 16983 7527 16989
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 8662 16980 8668 16992
rect 7515 16952 8668 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9582 16980 9588 16992
rect 9543 16952 9588 16980
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9824 16952 10241 16980
rect 9824 16940 9830 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10229 16943 10287 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 12342 16980 12348 16992
rect 12303 16952 12348 16980
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12492 16952 13001 16980
rect 12492 16940 12498 16952
rect 12989 16949 13001 16952
rect 13035 16949 13047 16983
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 12989 16943 13047 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15838 16980 15844 16992
rect 15799 16952 15844 16980
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 18874 16980 18880 16992
rect 17635 16952 18880 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 19334 16980 19340 16992
rect 19295 16952 19340 16980
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 19705 16983 19763 16989
rect 19705 16949 19717 16983
rect 19751 16980 19763 16983
rect 20070 16980 20076 16992
rect 19751 16952 20076 16980
rect 19751 16949 19763 16952
rect 19705 16943 19763 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 1104 16890 21436 16912
rect 1104 16838 4338 16890
rect 4390 16838 4402 16890
rect 4454 16838 4466 16890
rect 4518 16838 4530 16890
rect 4582 16838 4594 16890
rect 4646 16838 11116 16890
rect 11168 16838 11180 16890
rect 11232 16838 11244 16890
rect 11296 16838 11308 16890
rect 11360 16838 11372 16890
rect 11424 16838 17893 16890
rect 17945 16838 17957 16890
rect 18009 16838 18021 16890
rect 18073 16838 18085 16890
rect 18137 16838 18149 16890
rect 18201 16838 21436 16890
rect 1104 16816 21436 16838
rect 3605 16779 3663 16785
rect 3605 16745 3617 16779
rect 3651 16776 3663 16779
rect 4982 16776 4988 16788
rect 3651 16748 4988 16776
rect 3651 16745 3663 16748
rect 3605 16739 3663 16745
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 5224 16748 5273 16776
rect 5224 16736 5230 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 7101 16779 7159 16785
rect 7101 16745 7113 16779
rect 7147 16776 7159 16779
rect 7190 16776 7196 16788
rect 7147 16748 7196 16776
rect 7147 16745 7159 16748
rect 7101 16739 7159 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 9214 16776 9220 16788
rect 7432 16748 9220 16776
rect 7432 16736 7438 16748
rect 9214 16736 9220 16748
rect 9272 16776 9278 16788
rect 14182 16776 14188 16788
rect 9272 16748 14188 16776
rect 9272 16736 9278 16748
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14366 16776 14372 16788
rect 14327 16748 14372 16776
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 15565 16779 15623 16785
rect 15565 16776 15577 16779
rect 15344 16748 15577 16776
rect 15344 16736 15350 16748
rect 15565 16745 15577 16748
rect 15611 16745 15623 16779
rect 15565 16739 15623 16745
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 16114 16776 16120 16788
rect 16071 16748 16120 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17218 16776 17224 16788
rect 16816 16748 17224 16776
rect 16816 16736 16822 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19610 16776 19616 16788
rect 19475 16748 19616 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 3973 16711 4031 16717
rect 3973 16677 3985 16711
rect 4019 16677 4031 16711
rect 3973 16671 4031 16677
rect 1302 16532 1308 16584
rect 1360 16572 1366 16584
rect 2038 16572 2044 16584
rect 1360 16544 2044 16572
rect 1360 16532 1366 16544
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 2774 16572 2780 16584
rect 2547 16544 2780 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3292 16544 3801 16572
rect 3292 16532 3298 16544
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3988 16572 4016 16671
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 6880 16680 7297 16708
rect 6880 16668 6886 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 5092 16612 5304 16640
rect 4246 16572 4252 16584
rect 3988 16544 4252 16572
rect 3789 16535 3847 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16572 4491 16575
rect 4706 16572 4712 16584
rect 4479 16544 4712 16572
rect 4479 16541 4491 16544
rect 4433 16535 4491 16541
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 5092 16581 5120 16612
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16541 5135 16575
rect 5077 16535 5135 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5276 16572 5304 16612
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 7300 16640 7328 16671
rect 8846 16668 8852 16720
rect 8904 16708 8910 16720
rect 13722 16708 13728 16720
rect 8904 16680 13728 16708
rect 8904 16668 8910 16680
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 18046 16708 18052 16720
rect 14056 16680 18052 16708
rect 14056 16668 14062 16680
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 19702 16708 19708 16720
rect 18156 16680 19708 16708
rect 5408 16612 5453 16640
rect 7300 16612 7696 16640
rect 5408 16600 5414 16612
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 5276 16544 5917 16572
rect 5169 16535 5227 16541
rect 5905 16541 5917 16544
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 7006 16572 7012 16584
rect 6871 16544 7012 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 3605 16507 3663 16513
rect 3605 16504 3617 16507
rect 1872 16476 3617 16504
rect 1872 16445 1900 16476
rect 3605 16473 3617 16476
rect 3651 16473 3663 16507
rect 3605 16467 3663 16473
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 5184 16504 5212 16535
rect 3936 16476 5212 16504
rect 5920 16504 5948 16535
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16572 7251 16575
rect 7282 16572 7288 16584
rect 7239 16544 7288 16572
rect 7239 16541 7251 16544
rect 7193 16535 7251 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7524 16544 7573 16572
rect 7524 16532 7530 16544
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 7668 16572 7696 16612
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 10226 16640 10232 16652
rect 9364 16612 10232 16640
rect 9364 16600 9370 16612
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10410 16640 10416 16652
rect 10371 16612 10416 16640
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 12066 16640 12072 16652
rect 11532 16612 12072 16640
rect 10428 16572 10456 16600
rect 11532 16581 11560 16612
rect 12066 16600 12072 16612
rect 12124 16640 12130 16652
rect 12710 16640 12716 16652
rect 12124 16612 12716 16640
rect 12124 16600 12130 16612
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 14366 16640 14372 16652
rect 14139 16612 14372 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14366 16600 14372 16612
rect 14424 16640 14430 16652
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 14424 16612 14657 16640
rect 14424 16600 14430 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 14752 16612 16436 16640
rect 7668 16544 10456 16572
rect 11517 16575 11575 16581
rect 7561 16535 7619 16541
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 12897 16575 12955 16581
rect 12897 16572 12909 16575
rect 11756 16544 12909 16572
rect 11756 16532 11762 16544
rect 12897 16541 12909 16544
rect 12943 16572 12955 16575
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 12943 16544 13553 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 13541 16541 13553 16544
rect 13587 16572 13599 16575
rect 13630 16572 13636 16584
rect 13587 16544 13636 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 13630 16532 13636 16544
rect 13688 16572 13694 16584
rect 14274 16572 14280 16584
rect 13688 16544 14044 16572
rect 14235 16544 14280 16572
rect 13688 16532 13694 16544
rect 7374 16504 7380 16516
rect 5920 16476 7380 16504
rect 3936 16464 3942 16476
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 8110 16504 8116 16516
rect 7484 16476 8116 16504
rect 1857 16439 1915 16445
rect 1857 16405 1869 16439
rect 1903 16405 1915 16439
rect 2682 16436 2688 16448
rect 2643 16408 2688 16436
rect 1857 16399 1915 16405
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 4120 16408 4629 16436
rect 4120 16396 4126 16408
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 4890 16396 4896 16448
rect 4948 16436 4954 16448
rect 5718 16436 5724 16448
rect 4948 16408 5724 16436
rect 4948 16396 4954 16408
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16436 6055 16439
rect 7190 16436 7196 16448
rect 6043 16408 7196 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 7484 16445 7512 16476
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 9674 16464 9680 16516
rect 9732 16504 9738 16516
rect 13906 16504 13912 16516
rect 9732 16476 9904 16504
rect 9732 16464 9738 16476
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16405 7527 16439
rect 7469 16399 7527 16405
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 9769 16439 9827 16445
rect 9769 16436 9781 16439
rect 7708 16408 9781 16436
rect 7708 16396 7714 16408
rect 9769 16405 9781 16408
rect 9815 16405 9827 16439
rect 9876 16436 9904 16476
rect 12728 16476 13912 16504
rect 10137 16439 10195 16445
rect 10137 16436 10149 16439
rect 9876 16408 10149 16436
rect 9769 16399 9827 16405
rect 10137 16405 10149 16408
rect 10183 16405 10195 16439
rect 10137 16399 10195 16405
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10284 16408 10329 16436
rect 10284 16396 10290 16408
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11701 16439 11759 16445
rect 11701 16436 11713 16439
rect 11020 16408 11713 16436
rect 11020 16396 11026 16408
rect 11701 16405 11713 16408
rect 11747 16436 11759 16439
rect 11974 16436 11980 16448
rect 11747 16408 11980 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12728 16445 12756 16476
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 14016 16504 14044 16544
rect 14274 16532 14280 16544
rect 14332 16572 14338 16584
rect 14507 16575 14565 16581
rect 14507 16572 14519 16575
rect 14332 16544 14519 16572
rect 14332 16532 14338 16544
rect 14507 16541 14519 16544
rect 14553 16541 14565 16575
rect 14507 16535 14565 16541
rect 14752 16504 14780 16612
rect 16408 16584 16436 16612
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 17681 16643 17739 16649
rect 17681 16640 17693 16643
rect 16540 16612 17693 16640
rect 16540 16600 16546 16612
rect 17681 16609 17693 16612
rect 17727 16640 17739 16643
rect 18156 16640 18184 16680
rect 19702 16668 19708 16680
rect 19760 16668 19766 16720
rect 17727 16612 18184 16640
rect 18233 16643 18291 16649
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 18233 16609 18245 16643
rect 18279 16640 18291 16643
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 18279 16612 19901 16640
rect 18279 16609 18291 16612
rect 18233 16603 18291 16609
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20346 16640 20352 16652
rect 20119 16612 20352 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15436 16544 15577 16572
rect 15436 16532 15442 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 15930 16572 15936 16584
rect 15887 16544 15936 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 14016 16476 14780 16504
rect 14918 16464 14924 16516
rect 14976 16504 14982 16516
rect 15764 16504 15792 16535
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 14976 16476 15792 16504
rect 16132 16504 16160 16535
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16758 16572 16764 16584
rect 16448 16544 16764 16572
rect 16448 16532 16454 16544
rect 16758 16532 16764 16544
rect 16816 16572 16822 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16816 16544 16957 16572
rect 16816 16532 16822 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17034 16532 17040 16584
rect 17092 16572 17098 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17092 16544 17417 16572
rect 17092 16532 17098 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17552 16544 17597 16572
rect 17552 16532 17558 16544
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18417 16575 18475 16581
rect 18417 16572 18429 16575
rect 18104 16544 18429 16572
rect 18104 16532 18110 16544
rect 18417 16541 18429 16544
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 18564 16544 18705 16572
rect 18564 16532 18570 16544
rect 18693 16541 18705 16544
rect 18739 16572 18751 16575
rect 18782 16572 18788 16584
rect 18739 16544 18788 16572
rect 18739 16541 18751 16544
rect 18693 16535 18751 16541
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 19797 16575 19855 16581
rect 19797 16572 19809 16575
rect 19392 16544 19809 16572
rect 19392 16532 19398 16544
rect 19797 16541 19809 16544
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 17052 16504 17080 16532
rect 16132 16476 17080 16504
rect 14976 16464 14982 16476
rect 12713 16439 12771 16445
rect 12713 16405 12725 16439
rect 12759 16405 12771 16439
rect 12713 16399 12771 16405
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 15470 16436 15476 16448
rect 13403 16408 15476 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15764 16436 15792 16476
rect 16574 16436 16580 16448
rect 15764 16408 16580 16436
rect 16574 16396 16580 16408
rect 16632 16396 16638 16448
rect 16761 16439 16819 16445
rect 16761 16405 16773 16439
rect 16807 16436 16819 16439
rect 17126 16436 17132 16448
rect 16807 16408 17132 16436
rect 16807 16405 16819 16408
rect 16761 16399 16819 16405
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17678 16436 17684 16448
rect 17639 16408 17684 16436
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 18601 16439 18659 16445
rect 18601 16405 18613 16439
rect 18647 16436 18659 16439
rect 18874 16436 18880 16448
rect 18647 16408 18880 16436
rect 18647 16405 18659 16408
rect 18601 16399 18659 16405
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 1104 16346 21436 16368
rect 1104 16294 7727 16346
rect 7779 16294 7791 16346
rect 7843 16294 7855 16346
rect 7907 16294 7919 16346
rect 7971 16294 7983 16346
rect 8035 16294 14504 16346
rect 14556 16294 14568 16346
rect 14620 16294 14632 16346
rect 14684 16294 14696 16346
rect 14748 16294 14760 16346
rect 14812 16294 21436 16346
rect 1104 16272 21436 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1544 16204 1593 16232
rect 1544 16192 1550 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 3844 16204 4353 16232
rect 3844 16192 3850 16204
rect 4341 16201 4353 16204
rect 4387 16201 4399 16235
rect 4341 16195 4399 16201
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5077 16235 5135 16241
rect 5077 16232 5089 16235
rect 5040 16204 5089 16232
rect 5040 16192 5046 16204
rect 5077 16201 5089 16204
rect 5123 16201 5135 16235
rect 6270 16232 6276 16244
rect 5077 16195 5135 16201
rect 5184 16204 6276 16232
rect 1949 16167 2007 16173
rect 1949 16133 1961 16167
rect 1995 16164 2007 16167
rect 5184 16164 5212 16204
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 7098 16232 7104 16244
rect 7059 16204 7104 16232
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 10226 16192 10232 16244
rect 10284 16232 10290 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 10284 16204 12173 16232
rect 10284 16192 10290 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13320 16204 13461 16232
rect 13320 16192 13326 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 13449 16195 13507 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 17678 16232 17684 16244
rect 15528 16204 16804 16232
rect 17639 16204 17684 16232
rect 15528 16192 15534 16204
rect 1995 16136 5212 16164
rect 1995 16133 2007 16136
rect 1949 16127 2007 16133
rect 6362 16124 6368 16176
rect 6420 16164 6426 16176
rect 7193 16167 7251 16173
rect 7193 16164 7205 16167
rect 6420 16136 7205 16164
rect 6420 16124 6426 16136
rect 7193 16133 7205 16136
rect 7239 16133 7251 16167
rect 7193 16127 7251 16133
rect 8386 16124 8392 16176
rect 8444 16164 8450 16176
rect 10042 16164 10048 16176
rect 8444 16136 10048 16164
rect 8444 16124 8450 16136
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 11992 16136 12265 16164
rect 11992 16108 12020 16136
rect 12253 16133 12265 16136
rect 12299 16164 12311 16167
rect 12986 16164 12992 16176
rect 12299 16136 12992 16164
rect 12299 16133 12311 16136
rect 12253 16127 12311 16133
rect 12986 16124 12992 16136
rect 13044 16124 13050 16176
rect 14274 16124 14280 16176
rect 14332 16164 14338 16176
rect 14332 16136 14688 16164
rect 14332 16124 14338 16136
rect 3326 16096 3332 16108
rect 3287 16068 3332 16096
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3786 16096 3792 16108
rect 3651 16068 3792 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 4154 16096 4160 16108
rect 4115 16068 4160 16096
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 4847 16068 5488 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 2038 16028 2044 16040
rect 1999 16000 2044 16028
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2222 16028 2228 16040
rect 2183 16000 2228 16028
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3237 16031 3295 16037
rect 3237 16028 3249 16031
rect 2924 16000 3249 16028
rect 2924 15988 2930 16000
rect 3237 15997 3249 16000
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 15997 3755 16031
rect 5074 16028 5080 16040
rect 5035 16000 5080 16028
rect 3697 15991 3755 15997
rect 2240 15960 2268 15988
rect 3712 15960 3740 15991
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5460 16028 5488 16068
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5592 16068 5637 16096
rect 5592 16056 5598 16068
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5776 16068 5821 16096
rect 5776 16056 5782 16068
rect 7650 16056 7656 16108
rect 7708 16096 7714 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 7708 16068 10333 16096
rect 7708 16056 7714 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10468 16068 10517 16096
rect 10468 16056 10474 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 11974 16096 11980 16108
rect 11887 16068 11980 16096
rect 10505 16059 10563 16065
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 12802 16096 12808 16108
rect 12763 16068 12808 16096
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13814 16096 13820 16108
rect 13495 16068 13820 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14660 16105 14688 16136
rect 15010 16124 15016 16176
rect 15068 16164 15074 16176
rect 15068 16136 15976 16164
rect 15068 16124 15074 16136
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 14967 16068 15669 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 5810 16028 5816 16040
rect 5460 16000 5816 16028
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 6822 16028 6828 16040
rect 5920 16000 6828 16028
rect 4154 15960 4160 15972
rect 2240 15932 3648 15960
rect 3712 15932 4160 15960
rect 3050 15892 3056 15904
rect 3011 15864 3056 15892
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 3620 15892 3648 15932
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 4890 15960 4896 15972
rect 4803 15932 4896 15960
rect 4890 15920 4896 15932
rect 4948 15960 4954 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 4948 15932 5549 15960
rect 4948 15920 4954 15932
rect 5537 15929 5549 15932
rect 5583 15929 5595 15963
rect 5537 15923 5595 15929
rect 5920 15892 5948 16000
rect 6822 15988 6828 16000
rect 6880 16028 6886 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6880 16000 7297 16028
rect 6880 15988 6886 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 16028 10103 16031
rect 10778 16028 10784 16040
rect 10091 16000 10784 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10778 15988 10784 16000
rect 10836 16028 10842 16040
rect 11514 16028 11520 16040
rect 10836 16000 11520 16028
rect 10836 15988 10842 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 11790 16028 11796 16040
rect 11751 16000 11796 16028
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 12342 16028 12348 16040
rect 12303 16000 12348 16028
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 16028 13783 16031
rect 14568 16028 14596 16056
rect 13771 16000 14596 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 8260 15932 10149 15960
rect 8260 15920 8266 15932
rect 10137 15929 10149 15932
rect 10183 15960 10195 15963
rect 13541 15963 13599 15969
rect 10183 15932 13492 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 6730 15892 6736 15904
rect 3620 15864 5948 15892
rect 6691 15864 6736 15892
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 9858 15892 9864 15904
rect 9815 15864 9864 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10226 15892 10232 15904
rect 10100 15864 10232 15892
rect 10100 15852 10106 15864
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 12894 15892 12900 15904
rect 12855 15864 12900 15892
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 13464 15892 13492 15932
rect 13541 15929 13553 15963
rect 13587 15960 13599 15963
rect 13630 15960 13636 15972
rect 13587 15932 13636 15960
rect 13587 15929 13599 15932
rect 13541 15923 13599 15929
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 13740 15932 14964 15960
rect 13740 15892 13768 15932
rect 13464 15864 13768 15892
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 14090 15892 14096 15904
rect 13872 15864 14096 15892
rect 13872 15852 13878 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 14366 15892 14372 15904
rect 14327 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 14826 15892 14832 15904
rect 14787 15864 14832 15892
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 14936 15892 14964 15932
rect 15562 15920 15568 15972
rect 15620 15960 15626 15972
rect 15672 15960 15700 16059
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 15948 16105 15976 16136
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15804 16068 15853 16096
rect 15804 16056 15810 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 16132 16028 16160 16059
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16776 16096 16804 16204
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 19153 16167 19211 16173
rect 19153 16164 19165 16167
rect 17184 16136 19165 16164
rect 17184 16124 17190 16136
rect 19153 16133 19165 16136
rect 19199 16133 19211 16167
rect 19153 16127 19211 16133
rect 18598 16096 18604 16108
rect 16776 16068 18604 16096
rect 16669 16059 16727 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 19300 16068 20177 16096
rect 19300 16056 19306 16068
rect 20165 16065 20177 16068
rect 20211 16096 20223 16099
rect 20530 16096 20536 16108
rect 20211 16068 20536 16096
rect 20211 16065 20223 16068
rect 20165 16059 20223 16065
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 17034 16028 17040 16040
rect 16132 16000 17040 16028
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17644 16000 17785 16028
rect 17644 15988 17650 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 16761 15963 16819 15969
rect 16761 15960 16773 15963
rect 15620 15932 16773 15960
rect 15620 15920 15626 15932
rect 16761 15929 16773 15932
rect 16807 15929 16819 15963
rect 16761 15923 16819 15929
rect 17678 15920 17684 15972
rect 17736 15960 17742 15972
rect 17880 15960 17908 15991
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 18840 16000 19809 16028
rect 18840 15988 18846 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 20254 16028 20260 16040
rect 20215 16000 20260 16028
rect 19797 15991 19855 15997
rect 17736 15932 17908 15960
rect 17736 15920 17742 15932
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 19337 15963 19395 15969
rect 19337 15960 19349 15963
rect 19300 15932 19349 15960
rect 19300 15920 19306 15932
rect 19337 15929 19349 15932
rect 19383 15929 19395 15963
rect 19812 15960 19840 15991
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 20714 15960 20720 15972
rect 19812 15932 20720 15960
rect 19337 15923 19395 15929
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 15654 15892 15660 15904
rect 14936 15864 15660 15892
rect 15654 15852 15660 15864
rect 15712 15892 15718 15904
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 15712 15864 15761 15892
rect 15712 15852 15718 15864
rect 15749 15861 15761 15864
rect 15795 15892 15807 15895
rect 16206 15892 16212 15904
rect 15795 15864 16212 15892
rect 15795 15861 15807 15864
rect 15749 15855 15807 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 16724 15864 17325 15892
rect 16724 15852 16730 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 17313 15855 17371 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 1104 15802 21436 15824
rect 1104 15750 4338 15802
rect 4390 15750 4402 15802
rect 4454 15750 4466 15802
rect 4518 15750 4530 15802
rect 4582 15750 4594 15802
rect 4646 15750 11116 15802
rect 11168 15750 11180 15802
rect 11232 15750 11244 15802
rect 11296 15750 11308 15802
rect 11360 15750 11372 15802
rect 11424 15750 17893 15802
rect 17945 15750 17957 15802
rect 18009 15750 18021 15802
rect 18073 15750 18085 15802
rect 18137 15750 18149 15802
rect 18201 15750 21436 15802
rect 1104 15728 21436 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2096 15660 2697 15688
rect 2096 15648 2102 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 3786 15648 3792 15700
rect 3844 15688 3850 15700
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 3844 15660 5365 15688
rect 3844 15648 3850 15660
rect 5353 15657 5365 15660
rect 5399 15657 5411 15691
rect 5353 15651 5411 15657
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8536 15660 8953 15688
rect 8536 15648 8542 15660
rect 8941 15657 8953 15660
rect 8987 15688 8999 15691
rect 9030 15688 9036 15700
rect 8987 15660 9036 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 11974 15688 11980 15700
rect 9861 15651 9919 15657
rect 11164 15660 11980 15688
rect 1762 15580 1768 15632
rect 1820 15620 1826 15632
rect 3970 15620 3976 15632
rect 1820 15592 3976 15620
rect 1820 15580 1826 15592
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 5258 15620 5264 15632
rect 4816 15592 5264 15620
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 4816 15561 4844 15592
rect 5258 15580 5264 15592
rect 5316 15620 5322 15632
rect 5316 15592 5948 15620
rect 5316 15580 5322 15592
rect 3145 15555 3203 15561
rect 3145 15552 3157 15555
rect 2648 15524 3157 15552
rect 2648 15512 2654 15524
rect 3145 15521 3157 15524
rect 3191 15521 3203 15555
rect 3145 15515 3203 15521
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 4982 15512 4988 15564
rect 5040 15552 5046 15564
rect 5920 15561 5948 15592
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 10042 15620 10048 15632
rect 6604 15592 10048 15620
rect 6604 15580 6610 15592
rect 10042 15580 10048 15592
rect 10100 15580 10106 15632
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 5040 15524 5825 15552
rect 5040 15512 5046 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7156 15524 7481 15552
rect 7156 15512 7162 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 7469 15515 7527 15521
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 7616 15524 7665 15552
rect 7616 15512 7622 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 9398 15552 9404 15564
rect 9171 15524 9404 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 9398 15512 9404 15524
rect 9456 15552 9462 15564
rect 9582 15552 9588 15564
rect 9456 15524 9588 15552
rect 9456 15512 9462 15524
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10594 15552 10600 15564
rect 10367 15524 10600 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 2682 15484 2688 15496
rect 1719 15456 2688 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 2832 15456 2881 15484
rect 2832 15444 2838 15456
rect 2869 15453 2881 15456
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3237 15487 3295 15493
rect 3016 15456 3061 15484
rect 3016 15444 3022 15456
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 3252 15416 3280 15447
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 5776 15456 6561 15484
rect 5776 15444 5782 15456
rect 6549 15453 6561 15456
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 6641 15487 6699 15493
rect 6641 15453 6653 15487
rect 6687 15484 6699 15487
rect 7374 15484 7380 15496
rect 6687 15456 7380 15484
rect 6687 15453 6699 15456
rect 6641 15447 6699 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 9214 15484 9220 15496
rect 9175 15456 9220 15484
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9858 15484 9864 15496
rect 9819 15456 9864 15484
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 10008 15456 10057 15484
rect 10008 15444 10014 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 10137 15447 10195 15453
rect 2556 15388 3280 15416
rect 4525 15419 4583 15425
rect 2556 15376 2562 15388
rect 4525 15385 4537 15419
rect 4571 15416 4583 15419
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 4571 15388 7665 15416
rect 4571 15385 4583 15388
rect 4525 15379 4583 15385
rect 7653 15385 7665 15388
rect 7699 15385 7711 15419
rect 7653 15379 7711 15385
rect 8941 15419 8999 15425
rect 8941 15385 8953 15419
rect 8987 15385 8999 15419
rect 10152 15416 10180 15447
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 11164 15493 11192 15660
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 14608 15660 15945 15688
rect 14608 15648 14614 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 17034 15688 17040 15700
rect 16995 15660 17040 15688
rect 15933 15651 15991 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 17586 15688 17592 15700
rect 17547 15660 17592 15688
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 18601 15691 18659 15697
rect 18601 15657 18613 15691
rect 18647 15688 18659 15691
rect 18690 15688 18696 15700
rect 18647 15660 18696 15688
rect 18647 15657 18659 15660
rect 18601 15651 18659 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 11790 15620 11796 15632
rect 11256 15592 11796 15620
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 10778 15416 10784 15428
rect 10152 15388 10784 15416
rect 8941 15379 8999 15385
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 3292 15320 4169 15348
rect 3292 15308 3298 15320
rect 4157 15317 4169 15320
rect 4203 15317 4215 15351
rect 4157 15311 4215 15317
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 5718 15348 5724 15360
rect 4672 15320 4717 15348
rect 5679 15320 5724 15348
rect 4672 15308 4678 15320
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 8294 15348 8300 15360
rect 6604 15320 8300 15348
rect 6604 15308 6610 15320
rect 8294 15308 8300 15320
rect 8352 15348 8358 15360
rect 8956 15348 8984 15379
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11072 15416 11100 15447
rect 11256 15416 11284 15592
rect 11790 15580 11796 15592
rect 11848 15620 11854 15632
rect 12342 15620 12348 15632
rect 11848 15592 12348 15620
rect 11848 15580 11854 15592
rect 12342 15580 12348 15592
rect 12400 15620 12406 15632
rect 12437 15623 12495 15629
rect 12437 15620 12449 15623
rect 12400 15592 12449 15620
rect 12400 15580 12406 15592
rect 12437 15589 12449 15592
rect 12483 15620 12495 15623
rect 13081 15623 13139 15629
rect 13081 15620 13093 15623
rect 12483 15592 13093 15620
rect 12483 15589 12495 15592
rect 12437 15583 12495 15589
rect 13081 15589 13093 15592
rect 13127 15589 13139 15623
rect 13081 15583 13139 15589
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 12894 15552 12900 15564
rect 11379 15524 12900 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 11900 15493 11928 15524
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 14568 15552 14596 15648
rect 13311 15524 14596 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 16666 15552 16672 15564
rect 14884 15524 16672 15552
rect 14884 15512 14890 15524
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11348 15456 11437 15484
rect 11348 15428 11376 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12032 15456 12265 15484
rect 12032 15444 12038 15456
rect 12253 15453 12265 15456
rect 12299 15484 12311 15487
rect 12802 15484 12808 15496
rect 12299 15456 12808 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 13630 15484 13636 15496
rect 13219 15456 13636 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 14366 15484 14372 15496
rect 14327 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 15396 15493 15424 15524
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15453 15439 15487
rect 15562 15484 15568 15496
rect 15523 15456 15568 15484
rect 15381 15447 15439 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 16114 15484 16120 15496
rect 15795 15456 16120 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 16991 15456 17816 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 11072 15388 11284 15416
rect 11330 15376 11336 15428
rect 11388 15416 11394 15428
rect 12069 15419 12127 15425
rect 12069 15416 12081 15419
rect 11388 15388 12081 15416
rect 11388 15376 11394 15388
rect 12069 15385 12081 15388
rect 12115 15385 12127 15419
rect 12069 15379 12127 15385
rect 12161 15419 12219 15425
rect 12161 15385 12173 15419
rect 12207 15416 12219 15419
rect 12894 15416 12900 15428
rect 12207 15388 12296 15416
rect 12855 15388 12900 15416
rect 12207 15385 12219 15388
rect 12161 15379 12219 15385
rect 12268 15360 12296 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 14976 15388 15669 15416
rect 14976 15376 14982 15388
rect 15657 15385 15669 15388
rect 15703 15385 15715 15419
rect 17586 15416 17592 15428
rect 17547 15388 17592 15416
rect 15657 15379 15715 15385
rect 17586 15376 17592 15388
rect 17644 15376 17650 15428
rect 8352 15320 8984 15348
rect 8352 15308 8358 15320
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 9088 15320 9413 15348
rect 9088 15308 9094 15320
rect 9401 15317 9413 15320
rect 9447 15317 9459 15351
rect 9401 15311 9459 15317
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11882 15348 11888 15360
rect 10919 15320 11888 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12250 15308 12256 15360
rect 12308 15308 12314 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12584 15320 13001 15348
rect 12584 15308 12590 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 14274 15308 14280 15360
rect 14332 15348 14338 15360
rect 17788 15357 17816 15456
rect 17862 15444 17868 15496
rect 17920 15484 17926 15496
rect 18322 15484 18328 15496
rect 17920 15456 18328 15484
rect 17920 15444 17926 15456
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18874 15484 18880 15496
rect 18555 15456 18880 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19208 15456 19257 15484
rect 19208 15444 19214 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19886 15484 19892 15496
rect 19847 15456 19892 15484
rect 19245 15447 19303 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 14332 15320 14473 15348
rect 14332 15308 14338 15320
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14461 15311 14519 15317
rect 17773 15351 17831 15357
rect 17773 15317 17785 15351
rect 17819 15348 17831 15351
rect 18230 15348 18236 15360
rect 17819 15320 18236 15348
rect 17819 15317 17831 15320
rect 17773 15311 17831 15317
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 19334 15348 19340 15360
rect 19295 15320 19340 15348
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 1104 15258 21436 15280
rect 1104 15206 7727 15258
rect 7779 15206 7791 15258
rect 7843 15206 7855 15258
rect 7907 15206 7919 15258
rect 7971 15206 7983 15258
rect 8035 15206 14504 15258
rect 14556 15206 14568 15258
rect 14620 15206 14632 15258
rect 14684 15206 14696 15258
rect 14748 15206 14760 15258
rect 14812 15206 21436 15258
rect 1104 15184 21436 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2958 15144 2964 15156
rect 2179 15116 2964 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 4798 15144 4804 15156
rect 4663 15116 4804 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15144 5411 15147
rect 5718 15144 5724 15156
rect 5399 15116 5724 15144
rect 5399 15113 5411 15116
rect 5353 15107 5411 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7650 15144 7656 15156
rect 7607 15116 7656 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10686 15144 10692 15156
rect 10008 15116 10692 15144
rect 10008 15104 10014 15116
rect 10686 15104 10692 15116
rect 10744 15144 10750 15156
rect 12250 15144 12256 15156
rect 10744 15116 12256 15144
rect 10744 15104 10750 15116
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 16022 15144 16028 15156
rect 15620 15116 16028 15144
rect 15620 15104 15626 15116
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 20070 15144 20076 15156
rect 17552 15116 20076 15144
rect 17552 15104 17558 15116
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 20438 15144 20444 15156
rect 20211 15116 20444 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 3234 15076 3240 15088
rect 2976 15048 3240 15076
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2590 15008 2596 15020
rect 2087 14980 2596 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 2976 15017 3004 15048
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 4433 15079 4491 15085
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4890 15076 4896 15088
rect 4479 15048 4896 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4890 15036 4896 15048
rect 4948 15036 4954 15088
rect 5994 15076 6000 15088
rect 5552 15048 6000 15076
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 4982 15008 4988 15020
rect 4755 14980 4988 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5552 15017 5580 15048
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 7374 15036 7380 15088
rect 7432 15076 7438 15088
rect 7432 15048 7696 15076
rect 7432 15036 7438 15048
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5537 14971 5595 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 7668 15017 7696 15048
rect 9214 15036 9220 15088
rect 9272 15076 9278 15088
rect 10045 15079 10103 15085
rect 10045 15076 10057 15079
rect 9272 15048 10057 15076
rect 9272 15036 9278 15048
rect 10045 15045 10057 15048
rect 10091 15045 10103 15079
rect 10045 15039 10103 15045
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 10192 15048 10237 15076
rect 10192 15036 10198 15048
rect 10594 15036 10600 15088
rect 10652 15076 10658 15088
rect 10652 15048 12480 15076
rect 10652 15036 10658 15048
rect 12452 15020 12480 15048
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 12584 15048 12629 15076
rect 12584 15036 12590 15048
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 14976 15048 15976 15076
rect 14976 15036 14982 15048
rect 7653 15011 7711 15017
rect 5920 14980 6132 15008
rect 2866 14940 2872 14952
rect 2779 14912 2872 14940
rect 2866 14900 2872 14912
rect 2924 14940 2930 14952
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 2924 14912 3341 14940
rect 2924 14900 2930 14912
rect 3329 14909 3341 14912
rect 3375 14940 3387 14943
rect 5920 14940 5948 14980
rect 3375 14912 5948 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 4433 14875 4491 14881
rect 4433 14841 4445 14875
rect 4479 14872 4491 14875
rect 4614 14872 4620 14884
rect 4479 14844 4620 14872
rect 4479 14841 4491 14844
rect 4433 14835 4491 14841
rect 4614 14832 4620 14844
rect 4672 14832 4678 14884
rect 6104 14872 6132 14980
rect 7653 14977 7665 15011
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 10686 15008 10692 15020
rect 7800 14980 10088 15008
rect 10599 14980 10692 15008
rect 7800 14968 7806 14980
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6972 14912 7297 14940
rect 6972 14900 6978 14912
rect 7285 14909 7297 14912
rect 7331 14940 7343 14943
rect 8202 14940 8208 14952
rect 7331 14912 8208 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9950 14940 9956 14952
rect 9911 14912 9956 14940
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10060 14940 10088 14980
rect 10686 14968 10692 14980
rect 10744 15008 10750 15020
rect 11514 15008 11520 15020
rect 10744 14980 11520 15008
rect 10744 14968 10750 14980
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 12066 15008 12072 15020
rect 12027 14980 12072 15008
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 12434 14968 12440 15020
rect 12492 14968 12498 15020
rect 12618 15008 12624 15020
rect 12579 14980 12624 15008
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13446 15008 13452 15020
rect 13407 14980 13452 15008
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14093 15011 14151 15017
rect 14093 15008 14105 15011
rect 14056 14980 14105 15008
rect 14056 14968 14062 14980
rect 14093 14977 14105 14980
rect 14139 14977 14151 15011
rect 14093 14971 14151 14977
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14332 14980 14381 15008
rect 14332 14968 14338 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 15654 15008 15660 15020
rect 14875 14980 15660 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 12342 14949 12348 14952
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 10060 14912 11897 14940
rect 11885 14909 11897 14912
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 12328 14943 12348 14949
rect 12328 14909 12340 14943
rect 12328 14903 12348 14909
rect 12342 14900 12348 14903
rect 12400 14900 12406 14952
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 13044 14912 14473 14940
rect 13044 14900 13050 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14660 14940 14688 14971
rect 15654 14968 15660 14980
rect 15712 15008 15718 15020
rect 15948 15017 15976 15048
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 19702 15076 19708 15088
rect 17736 15048 19708 15076
rect 17736 15036 17742 15048
rect 19702 15036 19708 15048
rect 19760 15076 19766 15088
rect 20346 15076 20352 15088
rect 19760 15048 20352 15076
rect 19760 15036 19766 15048
rect 15749 15011 15807 15017
rect 15749 15008 15761 15011
rect 15712 14980 15761 15008
rect 15712 14968 15718 14980
rect 15749 14977 15761 14980
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 14977 15899 15011
rect 15841 14971 15899 14977
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 15856 14940 15884 14971
rect 16114 14968 16120 15020
rect 16172 15008 16178 15020
rect 16666 15008 16672 15020
rect 16172 14980 16265 15008
rect 16627 14980 16672 15008
rect 16172 14968 16178 14980
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 17862 15008 17868 15020
rect 17552 14980 17868 15008
rect 17552 14968 17558 14980
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 15008 18107 15011
rect 18230 15008 18236 15020
rect 18095 14980 18236 15008
rect 18095 14977 18107 14980
rect 18049 14971 18107 14977
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 14977 19119 15011
rect 19061 14971 19119 14977
rect 16022 14940 16028 14952
rect 14660 14912 16028 14940
rect 14461 14903 14519 14909
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 16132 14940 16160 14968
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16132 14912 16773 14940
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16761 14903 16819 14909
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 19076 14940 19104 14971
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19484 14980 20085 15008
rect 19484 14968 19490 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20272 14949 20300 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 16908 14912 19104 14940
rect 20257 14943 20315 14949
rect 16908 14900 16914 14912
rect 20257 14909 20269 14943
rect 20303 14909 20315 14943
rect 20257 14903 20315 14909
rect 7193 14875 7251 14881
rect 7193 14872 7205 14875
rect 6104 14844 7205 14872
rect 7193 14841 7205 14844
rect 7239 14872 7251 14875
rect 8110 14872 8116 14884
rect 7239 14844 8116 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 8110 14832 8116 14844
rect 8168 14832 8174 14884
rect 9585 14875 9643 14881
rect 9585 14841 9597 14875
rect 9631 14872 9643 14875
rect 11974 14872 11980 14884
rect 9631 14844 11980 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 16390 14832 16396 14884
rect 16448 14872 16454 14884
rect 17770 14872 17776 14884
rect 16448 14844 17776 14872
rect 16448 14832 16454 14844
rect 17770 14832 17776 14844
rect 17828 14872 17834 14884
rect 18322 14872 18328 14884
rect 17828 14844 18328 14872
rect 17828 14832 17834 14844
rect 18322 14832 18328 14844
rect 18380 14832 18386 14884
rect 19242 14872 19248 14884
rect 19203 14844 19248 14872
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2648 14776 2697 14804
rect 2648 14764 2654 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 5350 14804 5356 14816
rect 4856 14776 5356 14804
rect 4856 14764 4862 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5718 14804 5724 14816
rect 5679 14776 5724 14804
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 6917 14807 6975 14813
rect 6917 14804 6929 14807
rect 6880 14776 6929 14804
rect 6880 14764 6886 14776
rect 6917 14773 6929 14776
rect 6963 14773 6975 14807
rect 6917 14767 6975 14773
rect 7377 14807 7435 14813
rect 7377 14773 7389 14807
rect 7423 14804 7435 14807
rect 8386 14804 8392 14816
rect 7423 14776 8392 14804
rect 7423 14773 7435 14776
rect 7377 14767 7435 14773
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9674 14804 9680 14816
rect 8904 14776 9680 14804
rect 8904 14764 8910 14776
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10410 14804 10416 14816
rect 10192 14776 10416 14804
rect 10192 14764 10198 14776
rect 10410 14764 10416 14776
rect 10468 14804 10474 14816
rect 10781 14807 10839 14813
rect 10781 14804 10793 14807
rect 10468 14776 10793 14804
rect 10468 14764 10474 14776
rect 10781 14773 10793 14776
rect 10827 14773 10839 14807
rect 10781 14767 10839 14773
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13630 14804 13636 14816
rect 13587 14776 13636 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 15470 14804 15476 14816
rect 15431 14776 15476 14804
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17586 14804 17592 14816
rect 17184 14776 17592 14804
rect 17184 14764 17190 14776
rect 17586 14764 17592 14776
rect 17644 14804 17650 14816
rect 17865 14807 17923 14813
rect 17865 14804 17877 14807
rect 17644 14776 17877 14804
rect 17644 14764 17650 14776
rect 17865 14773 17877 14776
rect 17911 14773 17923 14807
rect 17865 14767 17923 14773
rect 19705 14807 19763 14813
rect 19705 14773 19717 14807
rect 19751 14804 19763 14807
rect 20438 14804 20444 14816
rect 19751 14776 20444 14804
rect 19751 14773 19763 14776
rect 19705 14767 19763 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 1104 14714 21436 14736
rect 1104 14662 4338 14714
rect 4390 14662 4402 14714
rect 4454 14662 4466 14714
rect 4518 14662 4530 14714
rect 4582 14662 4594 14714
rect 4646 14662 11116 14714
rect 11168 14662 11180 14714
rect 11232 14662 11244 14714
rect 11296 14662 11308 14714
rect 11360 14662 11372 14714
rect 11424 14662 17893 14714
rect 17945 14662 17957 14714
rect 18009 14662 18021 14714
rect 18073 14662 18085 14714
rect 18137 14662 18149 14714
rect 18201 14662 21436 14714
rect 1104 14640 21436 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 3234 14600 3240 14612
rect 2823 14572 3240 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4893 14603 4951 14609
rect 4893 14600 4905 14603
rect 4304 14572 4905 14600
rect 4304 14560 4310 14572
rect 4893 14569 4905 14572
rect 4939 14569 4951 14603
rect 4893 14563 4951 14569
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14532 2375 14535
rect 2406 14532 2412 14544
rect 2363 14504 2412 14532
rect 2363 14501 2375 14504
rect 2317 14495 2375 14501
rect 2406 14492 2412 14504
rect 2464 14532 2470 14544
rect 2464 14504 3832 14532
rect 2464 14492 2470 14504
rect 1762 14356 1768 14408
rect 1820 14396 1826 14408
rect 2498 14396 2504 14408
rect 1820 14368 2504 14396
rect 1820 14356 1826 14368
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2590 14356 2596 14408
rect 2648 14396 2654 14408
rect 2866 14396 2872 14408
rect 2648 14368 2693 14396
rect 2827 14368 2872 14396
rect 2648 14356 2654 14368
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3804 14405 3832 14504
rect 4908 14464 4936 14563
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 5132 14572 5273 14600
rect 5132 14560 5138 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5261 14563 5319 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6270 14560 6276 14612
rect 6328 14600 6334 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6328 14572 6929 14600
rect 6328 14560 6334 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 6917 14563 6975 14569
rect 7558 14560 7564 14612
rect 7616 14560 7622 14612
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9272 14572 9689 14600
rect 9272 14560 9278 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 10100 14572 10609 14600
rect 10100 14560 10106 14572
rect 10597 14569 10609 14572
rect 10643 14569 10655 14603
rect 10597 14563 10655 14569
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12124 14572 12449 14600
rect 12124 14560 12130 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 12437 14563 12495 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14553 14603 14611 14609
rect 14553 14600 14565 14603
rect 14332 14572 14565 14600
rect 14332 14560 14338 14572
rect 14553 14569 14565 14572
rect 14599 14569 14611 14603
rect 14553 14563 14611 14569
rect 16393 14603 16451 14609
rect 16393 14569 16405 14603
rect 16439 14600 16451 14603
rect 16850 14600 16856 14612
rect 16439 14572 16856 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17126 14600 17132 14612
rect 17087 14572 17132 14600
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17828 14572 17877 14600
rect 17828 14560 17834 14572
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 17865 14563 17923 14569
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 20714 14600 20720 14612
rect 20675 14572 20720 14600
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 7576 14532 7604 14560
rect 10778 14532 10784 14544
rect 7576 14504 7696 14532
rect 5166 14464 5172 14476
rect 4908 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 7190 14464 7196 14476
rect 5224 14436 5764 14464
rect 7151 14436 7196 14464
rect 5224 14424 5230 14436
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5350 14396 5356 14408
rect 5123 14368 5356 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 1670 14328 1676 14340
rect 1631 14300 1676 14328
rect 1670 14288 1676 14300
rect 1728 14288 1734 14340
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 4908 14328 4936 14359
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5736 14405 5764 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7432 14436 7573 14464
rect 7432 14424 7438 14436
rect 7561 14433 7573 14436
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14365 5779 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 5721 14359 5779 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7668 14405 7696 14504
rect 9646 14504 10784 14532
rect 9646 14464 9674 14504
rect 10778 14492 10784 14504
rect 10836 14532 10842 14544
rect 10965 14535 11023 14541
rect 10965 14532 10977 14535
rect 10836 14504 10977 14532
rect 10836 14492 10842 14504
rect 10965 14501 10977 14504
rect 11011 14501 11023 14535
rect 12897 14535 12955 14541
rect 12897 14532 12909 14535
rect 10965 14495 11023 14501
rect 11808 14504 12909 14532
rect 10686 14464 10692 14476
rect 7760 14436 9674 14464
rect 10060 14436 10692 14464
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 4982 14328 4988 14340
rect 1903 14300 4844 14328
rect 4908 14300 4988 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4816 14260 4844 14300
rect 4982 14288 4988 14300
rect 5040 14328 5046 14340
rect 5534 14328 5540 14340
rect 5040 14300 5540 14328
rect 5040 14288 5046 14300
rect 5534 14288 5540 14300
rect 5592 14328 5598 14340
rect 7760 14328 7788 14436
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9033 14399 9091 14405
rect 9033 14396 9045 14399
rect 8904 14368 9045 14396
rect 8904 14356 8910 14368
rect 9033 14365 9045 14368
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9306 14396 9312 14408
rect 9263 14368 9312 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 10060 14405 10088 14436
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10045 14399 10103 14405
rect 9916 14368 9961 14396
rect 9916 14356 9922 14368
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10594 14396 10600 14408
rect 10183 14368 10600 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 11808 14405 11836 14504
rect 12897 14501 12909 14504
rect 12943 14501 12955 14535
rect 12897 14495 12955 14501
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 15470 14532 15476 14544
rect 13219 14504 15476 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 18233 14535 18291 14541
rect 18233 14532 18245 14535
rect 17328 14504 18245 14532
rect 12066 14424 12072 14476
rect 12124 14424 12130 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 12912 14436 13369 14464
rect 11974 14405 11980 14408
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11941 14399 11980 14405
rect 11941 14365 11953 14399
rect 11941 14359 11980 14365
rect 11974 14356 11980 14359
rect 12032 14356 12038 14408
rect 12084 14396 12112 14424
rect 12277 14399 12335 14405
rect 12277 14396 12289 14399
rect 12084 14368 12289 14396
rect 12277 14365 12289 14368
rect 12323 14396 12335 14399
rect 12912 14396 12940 14436
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13504 14436 14688 14464
rect 13504 14424 13510 14436
rect 12323 14368 12940 14396
rect 13081 14399 13139 14405
rect 12323 14365 12335 14368
rect 12277 14359 12335 14365
rect 13081 14365 13093 14399
rect 13127 14365 13139 14399
rect 13262 14396 13268 14408
rect 13223 14368 13268 14396
rect 13081 14359 13139 14365
rect 5592 14300 7788 14328
rect 9125 14331 9183 14337
rect 5592 14288 5598 14300
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9171 14300 9996 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 8846 14260 8852 14272
rect 4816 14232 8852 14260
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 9968 14260 9996 14300
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 12066 14328 12072 14340
rect 11756 14300 12072 14328
rect 11756 14288 11762 14300
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14297 12219 14331
rect 13096 14328 13124 14359
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13538 14396 13544 14408
rect 13499 14368 13544 14396
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13688 14368 14289 14396
rect 13688 14356 13694 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14660 14405 14688 14436
rect 14734 14424 14740 14476
rect 14792 14464 14798 14476
rect 17328 14473 17356 14504
rect 18233 14501 18245 14504
rect 18279 14501 18291 14535
rect 18233 14495 18291 14501
rect 17313 14467 17371 14473
rect 17313 14464 17325 14467
rect 14792 14436 17325 14464
rect 14792 14424 14798 14436
rect 17313 14433 17325 14436
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 19392 14436 19901 14464
rect 19392 14424 19398 14436
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 14645 14399 14703 14405
rect 14424 14368 14469 14396
rect 14424 14356 14430 14368
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 16022 14396 16028 14408
rect 15151 14368 16028 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16114 14356 16120 14408
rect 16172 14396 16178 14408
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 16172 14368 16589 14396
rect 16172 14356 16178 14368
rect 16577 14365 16589 14368
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 17000 14368 17049 14396
rect 17000 14356 17006 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17552 14368 17877 14396
rect 17552 14356 17558 14368
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14396 18015 14399
rect 18230 14396 18236 14408
rect 18003 14368 18236 14396
rect 18003 14365 18015 14368
rect 17957 14359 18015 14365
rect 18230 14356 18236 14368
rect 18288 14396 18294 14408
rect 19610 14396 19616 14408
rect 18288 14368 18460 14396
rect 19571 14368 19616 14396
rect 18288 14356 18294 14368
rect 13998 14328 14004 14340
rect 13096 14300 14004 14328
rect 12161 14291 12219 14297
rect 10686 14260 10692 14272
rect 9916 14232 10692 14260
rect 9916 14220 9922 14232
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12176 14260 12204 14291
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 12250 14260 12256 14272
rect 11848 14232 12256 14260
rect 11848 14220 11854 14232
rect 12250 14220 12256 14232
rect 12308 14260 12314 14272
rect 13538 14260 13544 14272
rect 12308 14232 13544 14260
rect 12308 14220 12314 14232
rect 13538 14220 13544 14232
rect 13596 14260 13602 14272
rect 14274 14260 14280 14272
rect 13596 14232 14280 14260
rect 13596 14220 13602 14232
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15197 14263 15255 14269
rect 15197 14260 15209 14263
rect 14884 14232 15209 14260
rect 14884 14220 14890 14232
rect 15197 14229 15209 14232
rect 15243 14229 15255 14263
rect 15197 14223 15255 14229
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 17184 14232 17325 14260
rect 17184 14220 17190 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 18432 14260 18460 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 20070 14396 20076 14408
rect 19843 14368 20076 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20530 14396 20536 14408
rect 20180 14368 20536 14396
rect 18506 14288 18512 14340
rect 18564 14328 18570 14340
rect 20180 14328 20208 14368
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 18564 14300 20208 14328
rect 18564 14288 18570 14300
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 20349 14331 20407 14337
rect 20349 14328 20361 14331
rect 20312 14300 20361 14328
rect 20312 14288 20318 14300
rect 20349 14297 20361 14300
rect 20395 14297 20407 14331
rect 20349 14291 20407 14297
rect 21545 14263 21603 14269
rect 21545 14260 21557 14263
rect 18432 14232 21557 14260
rect 17313 14223 17371 14229
rect 21545 14229 21557 14232
rect 21591 14229 21603 14263
rect 21545 14223 21603 14229
rect 1104 14170 21436 14192
rect 1104 14118 7727 14170
rect 7779 14118 7791 14170
rect 7843 14118 7855 14170
rect 7907 14118 7919 14170
rect 7971 14118 7983 14170
rect 8035 14118 14504 14170
rect 14556 14118 14568 14170
rect 14620 14118 14632 14170
rect 14684 14118 14696 14170
rect 14748 14118 14760 14170
rect 14812 14118 21436 14170
rect 1104 14096 21436 14118
rect 3326 14056 3332 14068
rect 3239 14028 3332 14056
rect 3326 14016 3332 14028
rect 3384 14056 3390 14068
rect 3384 14028 4568 14056
rect 3384 14016 3390 14028
rect 2958 13988 2964 14000
rect 2608 13960 2964 13988
rect 1486 13920 1492 13932
rect 1447 13892 1492 13920
rect 1486 13880 1492 13892
rect 1544 13880 1550 13932
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 2332 13852 2360 13883
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 2464 13892 2509 13920
rect 2464 13880 2470 13892
rect 2608 13861 2636 13960
rect 2958 13948 2964 13960
rect 3016 13988 3022 14000
rect 3878 13988 3884 14000
rect 3016 13960 3884 13988
rect 3016 13948 3022 13960
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 4540 13997 4568 14028
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 5408 14028 5549 14056
rect 5408 14016 5414 14028
rect 5537 14025 5549 14028
rect 5583 14025 5595 14059
rect 5537 14019 5595 14025
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6696 14028 6837 14056
rect 6696 14016 6702 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7650 14056 7656 14068
rect 7515 14028 7656 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7650 14016 7656 14028
rect 7708 14056 7714 14068
rect 8202 14056 8208 14068
rect 7708 14028 8208 14056
rect 7708 14016 7714 14028
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 9950 14056 9956 14068
rect 9723 14028 9956 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 11882 14056 11888 14068
rect 11843 14028 11888 14056
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 14099 14059 14157 14065
rect 14099 14056 14111 14059
rect 13504 14028 14111 14056
rect 13504 14016 13510 14028
rect 14099 14025 14111 14028
rect 14145 14025 14157 14059
rect 14099 14019 14157 14025
rect 16022 14016 16028 14068
rect 16080 14056 16086 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16080 14028 16681 14056
rect 16080 14016 16086 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 16669 14019 16727 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 17368 14028 18061 14056
rect 17368 14016 17374 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 19794 14056 19800 14068
rect 18288 14028 19800 14056
rect 18288 14016 18294 14028
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 19978 14056 19984 14068
rect 19939 14028 19984 14056
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 20438 14056 20444 14068
rect 20211 14028 20444 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 4525 13991 4583 13997
rect 4525 13957 4537 13991
rect 4571 13988 4583 13991
rect 6733 13991 6791 13997
rect 6733 13988 6745 13991
rect 4571 13960 6745 13988
rect 4571 13957 4583 13960
rect 4525 13951 4583 13957
rect 6733 13957 6745 13960
rect 6779 13957 6791 13991
rect 6733 13951 6791 13957
rect 7190 13948 7196 14000
rect 7248 13988 7254 14000
rect 7248 13960 8064 13988
rect 7248 13948 7254 13960
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 3142 13920 3148 13932
rect 3103 13892 3148 13920
rect 2685 13883 2743 13889
rect 2593 13855 2651 13861
rect 2332 13824 2544 13852
rect 2516 13784 2544 13824
rect 2593 13821 2605 13855
rect 2639 13821 2651 13855
rect 2700 13852 2728 13883
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 4433 13923 4491 13929
rect 3476 13892 3521 13920
rect 3476 13880 3482 13892
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4479 13892 4660 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 2700 13824 3188 13852
rect 2593 13815 2651 13821
rect 2774 13784 2780 13796
rect 2516 13756 2780 13784
rect 2774 13744 2780 13756
rect 2832 13744 2838 13796
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 2130 13716 2136 13728
rect 2091 13688 2136 13716
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 3160 13725 3188 13824
rect 4154 13812 4160 13864
rect 4212 13812 4218 13864
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 4172 13784 4200 13812
rect 4632 13784 4660 13892
rect 4982 13880 4988 13932
rect 5040 13920 5046 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 5040 13892 5089 13920
rect 5040 13880 5046 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5442 13920 5448 13932
rect 5399 13892 5448 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 8036 13929 8064 13960
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 8168 13960 8213 13988
rect 8168 13948 8174 13960
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 11698 13988 11704 14000
rect 8904 13960 11704 13988
rect 8904 13948 8910 13960
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 11900 13988 11928 14016
rect 11808 13960 11928 13988
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7524 13892 7573 13920
rect 7524 13880 7530 13892
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 10134 13920 10140 13932
rect 10095 13892 10140 13920
rect 9861 13883 9919 13889
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5718 13852 5724 13864
rect 5307 13824 5724 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 6880 13824 7328 13852
rect 6880 13812 6886 13824
rect 5534 13784 5540 13796
rect 3292 13756 5540 13784
rect 3292 13744 3298 13756
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 6733 13787 6791 13793
rect 6733 13753 6745 13787
rect 6779 13784 6791 13787
rect 6779 13756 6868 13784
rect 6779 13753 6791 13756
rect 6733 13747 6791 13753
rect 3145 13719 3203 13725
rect 3145 13685 3157 13719
rect 3191 13716 3203 13719
rect 3694 13716 3700 13728
rect 3191 13688 3700 13716
rect 3191 13685 3203 13688
rect 3145 13679 3203 13685
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 6840 13716 6868 13756
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7300 13793 7328 13824
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9876 13852 9904 13883
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10594 13920 10600 13932
rect 10555 13892 10600 13920
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 10744 13892 10789 13920
rect 10744 13880 10750 13892
rect 10410 13852 10416 13864
rect 8352 13824 10416 13852
rect 8352 13812 8358 13824
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10836 13824 10885 13852
rect 10836 13812 10842 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 11808 13852 11836 13960
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12250 13988 12256 14000
rect 12032 13960 12256 13988
rect 12032 13948 12038 13960
rect 12250 13948 12256 13960
rect 12308 13988 12314 14000
rect 12805 13991 12863 13997
rect 12805 13988 12817 13991
rect 12308 13960 12817 13988
rect 12308 13948 12314 13960
rect 12805 13957 12817 13960
rect 12851 13957 12863 13991
rect 14182 13988 14188 14000
rect 14095 13960 14188 13988
rect 12805 13951 12863 13957
rect 14182 13948 14188 13960
rect 14240 13988 14246 14000
rect 14240 13960 14964 13988
rect 14240 13948 14246 13960
rect 11882 13923 11940 13929
rect 11882 13889 11894 13923
rect 11928 13920 11940 13923
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 11928 13892 12357 13920
rect 11928 13889 11940 13892
rect 11882 13883 11940 13889
rect 12345 13889 12357 13892
rect 12391 13920 12403 13923
rect 12894 13920 12900 13932
rect 12391 13892 12900 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13920 13047 13923
rect 13998 13920 14004 13932
rect 13035 13892 13308 13920
rect 13911 13892 14004 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 11808 13824 12265 13852
rect 10873 13815 10931 13821
rect 12253 13821 12265 13824
rect 12299 13821 12311 13855
rect 13173 13855 13231 13861
rect 13173 13852 13185 13855
rect 12253 13815 12311 13821
rect 12452 13824 13185 13852
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 6972 13756 7205 13784
rect 6972 13744 6978 13756
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 7285 13787 7343 13793
rect 7285 13753 7297 13787
rect 7331 13784 7343 13787
rect 8386 13784 8392 13796
rect 7331 13756 8392 13784
rect 7331 13753 7343 13756
rect 7285 13747 7343 13753
rect 8386 13744 8392 13756
rect 8444 13744 8450 13796
rect 10045 13787 10103 13793
rect 10045 13753 10057 13787
rect 10091 13784 10103 13787
rect 10962 13784 10968 13796
rect 10091 13756 10968 13784
rect 10091 13753 10103 13756
rect 10045 13747 10103 13753
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 11974 13784 11980 13796
rect 11664 13756 11980 13784
rect 11664 13744 11670 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 12452 13784 12480 13824
rect 13173 13821 13185 13824
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 12400 13756 12480 13784
rect 12400 13744 12406 13756
rect 7101 13719 7159 13725
rect 7101 13716 7113 13719
rect 6840 13688 7113 13716
rect 7101 13685 7113 13688
rect 7147 13685 7159 13719
rect 7101 13679 7159 13685
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9398 13716 9404 13728
rect 9088 13688 9404 13716
rect 9088 13676 9094 13688
rect 9398 13676 9404 13688
rect 9456 13676 9462 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9950 13716 9956 13728
rect 9640 13688 9956 13716
rect 9640 13676 9646 13688
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10778 13716 10784 13728
rect 10739 13688 10784 13716
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 13280 13716 13308 13892
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 14323 13892 14749 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 14737 13889 14749 13892
rect 14783 13920 14795 13923
rect 14826 13920 14832 13932
rect 14783 13892 14832 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 14936 13929 14964 13960
rect 18598 13948 18604 14000
rect 18656 13988 18662 14000
rect 18656 13960 19196 13988
rect 18656 13948 18662 13960
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15746 13920 15752 13932
rect 15252 13892 15752 13920
rect 15252 13880 15258 13892
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 17034 13920 17040 13932
rect 16995 13892 17040 13920
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17678 13920 17684 13932
rect 17328 13892 17684 13920
rect 14016 13852 14044 13880
rect 17328 13861 17356 13892
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 19168 13929 19196 13960
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19702 13988 19708 14000
rect 19300 13960 19708 13988
rect 19300 13948 19306 13960
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18340 13920 18460 13926
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 17911 13898 18889 13920
rect 17911 13892 18368 13898
rect 18432 13892 18889 13898
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 17313 13855 17371 13861
rect 14016 13824 14780 13852
rect 13998 13744 14004 13796
rect 14056 13784 14062 13796
rect 14752 13793 14780 13824
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13821 18015 13855
rect 18138 13852 18144 13864
rect 18099 13824 18144 13852
rect 17957 13815 18015 13821
rect 14737 13787 14795 13793
rect 14056 13756 14688 13784
rect 14056 13744 14062 13756
rect 12124 13688 13308 13716
rect 14660 13716 14688 13756
rect 14737 13753 14749 13787
rect 14783 13753 14795 13787
rect 14737 13747 14795 13753
rect 14844 13756 17264 13784
rect 14844 13716 14872 13756
rect 14660 13688 14872 13716
rect 17236 13716 17264 13756
rect 17678 13744 17684 13796
rect 17736 13784 17742 13796
rect 17972 13784 18000 13815
rect 18138 13812 18144 13824
rect 18196 13812 18202 13864
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18380 13824 18429 13852
rect 18380 13812 18386 13824
rect 18417 13821 18429 13824
rect 18463 13821 18475 13855
rect 18417 13815 18475 13821
rect 19076 13852 19104 13883
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19392 13892 19441 13920
rect 19392 13880 19398 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19886 13920 19892 13932
rect 19429 13883 19487 13889
rect 19536 13892 19892 13920
rect 19536 13852 19564 13892
rect 19886 13880 19892 13892
rect 19944 13920 19950 13932
rect 20162 13920 20168 13932
rect 19944 13892 20168 13920
rect 19944 13880 19950 13892
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20530 13920 20536 13932
rect 20491 13892 20536 13920
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 19076 13824 19564 13852
rect 19076 13784 19104 13824
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20404 13824 20637 13852
rect 20404 13812 20410 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 17736 13756 19104 13784
rect 19245 13787 19303 13793
rect 17736 13744 17742 13756
rect 19245 13753 19257 13787
rect 19291 13784 19303 13787
rect 19518 13784 19524 13796
rect 19291 13756 19524 13784
rect 19291 13753 19303 13756
rect 19245 13747 19303 13753
rect 19518 13744 19524 13756
rect 19576 13744 19582 13796
rect 18230 13716 18236 13728
rect 17236 13688 18236 13716
rect 12124 13676 12130 13688
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18325 13719 18383 13725
rect 18325 13685 18337 13719
rect 18371 13716 18383 13719
rect 18506 13716 18512 13728
rect 18371 13688 18512 13716
rect 18371 13685 18383 13688
rect 18325 13679 18383 13685
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 19337 13719 19395 13725
rect 19337 13685 19349 13719
rect 19383 13716 19395 13719
rect 19426 13716 19432 13728
rect 19383 13688 19432 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 19426 13676 19432 13688
rect 19484 13716 19490 13728
rect 19794 13716 19800 13728
rect 19484 13688 19800 13716
rect 19484 13676 19490 13688
rect 19794 13676 19800 13688
rect 19852 13676 19858 13728
rect 1104 13626 21436 13648
rect 1104 13574 4338 13626
rect 4390 13574 4402 13626
rect 4454 13574 4466 13626
rect 4518 13574 4530 13626
rect 4582 13574 4594 13626
rect 4646 13574 11116 13626
rect 11168 13574 11180 13626
rect 11232 13574 11244 13626
rect 11296 13574 11308 13626
rect 11360 13574 11372 13626
rect 11424 13574 17893 13626
rect 17945 13574 17957 13626
rect 18009 13574 18021 13626
rect 18073 13574 18085 13626
rect 18137 13574 18149 13626
rect 18201 13574 21436 13626
rect 1104 13552 21436 13574
rect 2866 13512 2872 13524
rect 2779 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13512 2930 13524
rect 3142 13512 3148 13524
rect 2924 13484 3148 13512
rect 2924 13472 2930 13484
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 3476 13484 3893 13512
rect 3476 13472 3482 13484
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 3881 13475 3939 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 9306 13512 9312 13524
rect 9232 13484 9312 13512
rect 2130 13376 2136 13388
rect 2091 13348 2136 13376
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 3436 13376 3464 13472
rect 6454 13404 6460 13456
rect 6512 13444 6518 13456
rect 7650 13444 7656 13456
rect 6512 13416 7656 13444
rect 6512 13404 6518 13416
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 9232 13444 9260 13484
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10100 13484 11192 13512
rect 10100 13472 10106 13484
rect 8628 13416 9260 13444
rect 8628 13404 8634 13416
rect 5074 13376 5080 13388
rect 2280 13348 2325 13376
rect 2884 13348 3464 13376
rect 4724 13348 5080 13376
rect 2280 13336 2286 13348
rect 2884 13317 2912 13348
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3326 13308 3332 13320
rect 3099 13280 3332 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3418 13268 3424 13320
rect 3476 13308 3482 13320
rect 3786 13308 3792 13320
rect 3476 13280 3792 13308
rect 3476 13268 3482 13280
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 4724 13317 4752 13348
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 7101 13379 7159 13385
rect 5592 13348 6868 13376
rect 5592 13336 5598 13348
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 6638 13308 6644 13320
rect 4939 13280 5580 13308
rect 6599 13280 6644 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 2041 13243 2099 13249
rect 2041 13209 2053 13243
rect 2087 13240 2099 13243
rect 5353 13243 5411 13249
rect 2087 13212 4936 13240
rect 2087 13209 2099 13212
rect 2041 13203 2099 13209
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 2314 13172 2320 13184
rect 1719 13144 2320 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2682 13132 2688 13184
rect 2740 13172 2746 13184
rect 4614 13172 4620 13184
rect 2740 13144 4620 13172
rect 2740 13132 2746 13144
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4798 13172 4804 13184
rect 4759 13144 4804 13172
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 4908 13172 4936 13212
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 5442 13240 5448 13252
rect 5399 13212 5448 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 5552 13249 5580 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6840 13317 6868 13348
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7558 13376 7564 13388
rect 7147 13348 7564 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7558 13336 7564 13348
rect 7616 13376 7622 13388
rect 8110 13376 8116 13388
rect 7616 13348 8116 13376
rect 7616 13336 7622 13348
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8904 13348 9045 13376
rect 8904 13336 8910 13348
rect 9033 13345 9045 13348
rect 9079 13376 9091 13379
rect 9122 13376 9128 13388
rect 9079 13348 9128 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9232 13385 9260 13416
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 10134 13444 10140 13456
rect 9456 13416 10140 13444
rect 9456 13404 9462 13416
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 10226 13404 10232 13456
rect 10284 13444 10290 13456
rect 10284 13416 10548 13444
rect 10284 13404 10290 13416
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13345 9275 13379
rect 9217 13339 9275 13345
rect 9309 13379 9367 13385
rect 9309 13345 9321 13379
rect 9355 13376 9367 13379
rect 10042 13376 10048 13388
rect 9355 13348 10048 13376
rect 9355 13345 9367 13348
rect 9309 13339 9367 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10520 13385 10548 13416
rect 10778 13404 10784 13456
rect 10836 13404 10842 13456
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7466 13308 7472 13320
rect 7239 13280 7472 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 5537 13243 5595 13249
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 5810 13240 5816 13252
rect 5583 13212 5816 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 6641 13175 6699 13181
rect 6641 13172 6653 13175
rect 4908 13144 6653 13172
rect 6641 13141 6653 13144
rect 6687 13141 6699 13175
rect 6840 13172 6868 13271
rect 6932 13240 6960 13271
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 9490 13308 9496 13320
rect 8444 13280 9496 13308
rect 8444 13268 8450 13280
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10796 13308 10824 13404
rect 11164 13317 11192 13484
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 12342 13512 12348 13524
rect 11848 13484 12348 13512
rect 11848 13472 11854 13484
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12437 13515 12495 13521
rect 12437 13481 12449 13515
rect 12483 13512 12495 13515
rect 12894 13512 12900 13524
rect 12483 13484 12900 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 14182 13512 14188 13524
rect 14143 13484 14188 13512
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 14918 13512 14924 13524
rect 14879 13484 14924 13512
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 15933 13515 15991 13521
rect 15933 13481 15945 13515
rect 15979 13481 15991 13515
rect 15933 13475 15991 13481
rect 16945 13515 17003 13521
rect 16945 13481 16957 13515
rect 16991 13512 17003 13515
rect 17494 13512 17500 13524
rect 16991 13484 17500 13512
rect 16991 13481 17003 13484
rect 16945 13475 17003 13481
rect 15197 13447 15255 13453
rect 15197 13413 15209 13447
rect 15243 13444 15255 13447
rect 15948 13444 15976 13475
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17773 13515 17831 13521
rect 17773 13481 17785 13515
rect 17819 13512 17831 13515
rect 19702 13512 19708 13524
rect 17819 13484 19708 13512
rect 17819 13481 17831 13484
rect 17773 13475 17831 13481
rect 19702 13472 19708 13484
rect 19760 13512 19766 13524
rect 20530 13512 20536 13524
rect 19760 13484 20536 13512
rect 19760 13472 19766 13484
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 17129 13447 17187 13453
rect 17129 13444 17141 13447
rect 15243 13416 15792 13444
rect 15948 13416 17141 13444
rect 15243 13413 15255 13416
rect 15197 13407 15255 13413
rect 11790 13376 11796 13388
rect 11751 13348 11796 13376
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 15764 13385 15792 13416
rect 17129 13413 17141 13416
rect 17175 13413 17187 13447
rect 17129 13407 17187 13413
rect 18230 13404 18236 13456
rect 18288 13444 18294 13456
rect 19245 13447 19303 13453
rect 19245 13444 19257 13447
rect 18288 13416 19257 13444
rect 18288 13404 18294 13416
rect 19245 13413 19257 13416
rect 19291 13413 19303 13447
rect 20438 13444 20444 13456
rect 19245 13407 19303 13413
rect 19444 13416 20444 13444
rect 14829 13379 14887 13385
rect 14829 13376 14841 13379
rect 12176 13348 14841 13376
rect 10459 13280 10824 13308
rect 11149 13311 11207 13317
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 11149 13277 11161 13311
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12176 13317 12204 13348
rect 14829 13345 14841 13348
rect 14875 13345 14887 13379
rect 14829 13339 14887 13345
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 16574 13376 16580 13388
rect 16172 13348 16252 13376
rect 16487 13348 16580 13376
rect 16172 13336 16178 13348
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 12124 13280 12173 13308
rect 12124 13268 12130 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 14093 13311 14151 13317
rect 12308 13280 12401 13308
rect 12308 13268 12314 13280
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 7282 13240 7288 13252
rect 6932 13212 7288 13240
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 11256 13240 11284 13268
rect 9968 13212 11284 13240
rect 8846 13172 8852 13184
rect 6840 13144 8852 13172
rect 6641 13135 6699 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 9030 13172 9036 13184
rect 8991 13144 9036 13172
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9214 13172 9220 13184
rect 9171 13144 9220 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9968 13181 9996 13212
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 12268 13240 12296 13268
rect 11480 13212 12296 13240
rect 11480 13200 11486 13212
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 13998 13240 14004 13252
rect 12400 13212 14004 13240
rect 12400 13200 12406 13212
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14108 13240 14136 13271
rect 14274 13268 14280 13320
rect 14332 13308 14338 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14332 13280 14749 13308
rect 14332 13268 14338 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15470 13308 15476 13320
rect 15059 13280 15476 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 14366 13240 14372 13252
rect 14108 13212 14372 13240
rect 14366 13200 14372 13212
rect 14424 13240 14430 13252
rect 15028 13240 15056 13271
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 14424 13212 15056 13240
rect 15657 13243 15715 13249
rect 14424 13200 14430 13212
rect 15657 13209 15669 13243
rect 15703 13240 15715 13243
rect 15838 13240 15844 13252
rect 15703 13212 15844 13240
rect 15703 13209 15715 13212
rect 15657 13203 15715 13209
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 10284 13144 10333 13172
rect 10284 13132 10290 13144
rect 10321 13141 10333 13144
rect 10367 13141 10379 13175
rect 10321 13135 10379 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 10744 13144 11253 13172
rect 10744 13132 10750 13144
rect 11241 13141 11253 13144
rect 11287 13141 11299 13175
rect 11241 13135 11299 13141
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 15948 13172 15976 13271
rect 16224 13184 16252 13348
rect 16574 13336 16580 13348
rect 16632 13376 16638 13388
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 16632 13348 16773 13376
rect 16632 13336 16638 13348
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 16908 13348 18705 13376
rect 16908 13336 16914 13348
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17126 13308 17132 13320
rect 16991 13280 17132 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18046 13308 18052 13320
rect 18003 13280 18052 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 17678 13240 17684 13252
rect 16715 13212 17684 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 17788 13240 17816 13271
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 19444 13308 19472 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 20622 13376 20628 13388
rect 19935 13348 20628 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 18340 13280 19472 13308
rect 18340 13240 18368 13280
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19576 13280 19625 13308
rect 19576 13268 19582 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 18506 13240 18512 13252
rect 17788 13212 18368 13240
rect 18467 13212 18512 13240
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18598 13200 18604 13252
rect 18656 13240 18662 13252
rect 20533 13243 20591 13249
rect 18656 13212 19840 13240
rect 18656 13200 18662 13212
rect 16114 13172 16120 13184
rect 12676 13144 15976 13172
rect 16075 13144 16120 13172
rect 12676 13132 12682 13144
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16206 13132 16212 13184
rect 16264 13132 16270 13184
rect 16577 13175 16635 13181
rect 16577 13141 16589 13175
rect 16623 13172 16635 13175
rect 16850 13172 16856 13184
rect 16623 13144 16856 13172
rect 16623 13141 16635 13144
rect 16577 13135 16635 13141
rect 16850 13132 16856 13144
rect 16908 13132 16914 13184
rect 17696 13172 17724 13200
rect 18046 13172 18052 13184
rect 17696 13144 18052 13172
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19705 13175 19763 13181
rect 19705 13172 19717 13175
rect 19484 13144 19717 13172
rect 19484 13132 19490 13144
rect 19705 13141 19717 13144
rect 19751 13141 19763 13175
rect 19812 13172 19840 13212
rect 20533 13209 20545 13243
rect 20579 13240 20591 13243
rect 20714 13240 20720 13252
rect 20579 13212 20720 13240
rect 20579 13209 20591 13212
rect 20533 13203 20591 13209
rect 20714 13200 20720 13212
rect 20772 13200 20778 13252
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 19812 13144 20637 13172
rect 19705 13135 19763 13141
rect 20625 13141 20637 13144
rect 20671 13141 20683 13175
rect 20625 13135 20683 13141
rect 1104 13082 21436 13104
rect 1104 13030 7727 13082
rect 7779 13030 7791 13082
rect 7843 13030 7855 13082
rect 7907 13030 7919 13082
rect 7971 13030 7983 13082
rect 8035 13030 14504 13082
rect 14556 13030 14568 13082
rect 14620 13030 14632 13082
rect 14684 13030 14696 13082
rect 14748 13030 14760 13082
rect 14812 13030 21436 13082
rect 1104 13008 21436 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 6546 12968 6552 12980
rect 1995 12940 6552 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 9766 12968 9772 12980
rect 6840 12940 9772 12968
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3786 12900 3792 12912
rect 2832 12872 3792 12900
rect 2832 12860 2838 12872
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 5261 12903 5319 12909
rect 5261 12869 5273 12903
rect 5307 12900 5319 12903
rect 5810 12900 5816 12912
rect 5307 12872 5816 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 1854 12832 1860 12844
rect 1815 12804 1860 12832
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 2866 12832 2872 12844
rect 2827 12804 2872 12832
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3234 12832 3240 12844
rect 3016 12804 3061 12832
rect 3195 12804 3240 12832
rect 3016 12792 3022 12804
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3694 12832 3700 12844
rect 3655 12804 3700 12832
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4856 12804 5089 12832
rect 4856 12792 4862 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 3142 12764 3148 12776
rect 3055 12736 3148 12764
rect 3142 12724 3148 12736
rect 3200 12764 3206 12776
rect 3418 12764 3424 12776
rect 3200 12736 3424 12764
rect 3200 12724 3206 12736
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 5092 12764 5120 12795
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 5224 12804 5365 12832
rect 5224 12792 5230 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 6840 12841 6868 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10226 12968 10232 12980
rect 10187 12940 10232 12968
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10468 12940 10824 12968
rect 10468 12928 10474 12940
rect 7466 12900 7472 12912
rect 7427 12872 7472 12900
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 9122 12860 9128 12912
rect 9180 12900 9186 12912
rect 10686 12900 10692 12912
rect 9180 12872 9444 12900
rect 9180 12860 9186 12872
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 5500 12804 6837 12832
rect 5500 12792 5506 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 7650 12832 7656 12844
rect 7611 12804 7656 12832
rect 6825 12795 6883 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 8846 12832 8852 12844
rect 7791 12804 8852 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9416 12841 9444 12872
rect 9784 12872 10692 12900
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 9088 12804 9229 12832
rect 9088 12792 9094 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9582 12832 9588 12844
rect 9539 12804 9588 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 9784 12841 9812 12872
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 10796 12900 10824 12940
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11756 12940 11989 12968
rect 11756 12928 11762 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 13265 12971 13323 12977
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 14090 12968 14096 12980
rect 13311 12940 14096 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14645 12971 14703 12977
rect 14645 12937 14657 12971
rect 14691 12968 14703 12971
rect 15010 12968 15016 12980
rect 14691 12940 15016 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 17034 12968 17040 12980
rect 16715 12940 17040 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19613 12971 19671 12977
rect 19613 12937 19625 12971
rect 19659 12968 19671 12971
rect 19978 12968 19984 12980
rect 19659 12940 19984 12968
rect 19659 12937 19671 12940
rect 19613 12931 19671 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 11790 12900 11796 12912
rect 10796 12872 11796 12900
rect 11790 12860 11796 12872
rect 11848 12900 11854 12912
rect 11848 12872 16896 12900
rect 11848 12860 11854 12872
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 9769 12795 9827 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 10612 12804 11897 12832
rect 5534 12764 5540 12776
rect 5092 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6086 12764 6092 12776
rect 5684 12736 6092 12764
rect 5684 12724 5690 12736
rect 6086 12724 6092 12736
rect 6144 12764 6150 12776
rect 7466 12764 7472 12776
rect 6144 12736 7472 12764
rect 6144 12724 6150 12736
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 10612 12764 10640 12804
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13998 12832 14004 12844
rect 13219 12804 14004 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 14240 12804 14289 12832
rect 14240 12792 14246 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14734 12832 14740 12844
rect 14695 12804 14740 12832
rect 14277 12795 14335 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 16868 12841 16896 12872
rect 17402 12860 17408 12912
rect 17460 12900 17466 12912
rect 20162 12900 20168 12912
rect 17460 12872 20168 12900
rect 17460 12860 17466 12872
rect 20162 12860 20168 12872
rect 20220 12900 20226 12912
rect 20220 12872 20576 12900
rect 20220 12860 20226 12872
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16853 12835 16911 12841
rect 15979 12804 16068 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 9355 12736 10640 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 12161 12767 12219 12773
rect 10744 12736 10789 12764
rect 10744 12724 10750 12736
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12802 12764 12808 12776
rect 12207 12736 12808 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12802 12724 12808 12736
rect 12860 12764 12866 12776
rect 13262 12764 13268 12776
rect 12860 12736 13268 12764
rect 12860 12724 12866 12736
rect 13262 12724 13268 12736
rect 13320 12764 13326 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 13320 12736 13369 12764
rect 13320 12724 13326 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 13357 12727 13415 12733
rect 13464 12736 14473 12764
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 4672 12668 9444 12696
rect 4672 12656 4678 12668
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 6917 12631 6975 12637
rect 6917 12628 6929 12631
rect 6880 12600 6929 12628
rect 6880 12588 6886 12600
rect 6917 12597 6929 12600
rect 6963 12597 6975 12631
rect 6917 12591 6975 12597
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7466 12628 7472 12640
rect 7248 12600 7472 12628
rect 7248 12588 7254 12600
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7929 12631 7987 12637
rect 7929 12597 7941 12631
rect 7975 12628 7987 12631
rect 9122 12628 9128 12640
rect 7975 12600 9128 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9416 12628 9444 12668
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 9548 12668 9689 12696
rect 9548 12656 9554 12668
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 13464 12696 13492 12736
rect 14461 12733 14473 12736
rect 14507 12764 14519 12767
rect 15194 12764 15200 12776
rect 14507 12736 15200 12764
rect 14507 12733 14519 12736
rect 14461 12727 14519 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 16040 12764 16068 12804
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17368 12804 17601 12832
rect 17368 12792 17374 12804
rect 17589 12801 17601 12804
rect 17635 12832 17647 12835
rect 17770 12832 17776 12844
rect 17635 12804 17776 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18380 12804 18613 12832
rect 18380 12792 18386 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 19150 12792 19156 12844
rect 19208 12832 19214 12844
rect 19610 12835 19668 12841
rect 19610 12832 19622 12835
rect 19208 12804 19622 12832
rect 19208 12792 19214 12804
rect 19610 12801 19622 12804
rect 19656 12832 19668 12835
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19656 12804 20085 12832
rect 19656 12801 19668 12804
rect 19610 12795 19668 12801
rect 20073 12801 20085 12804
rect 20119 12832 20131 12835
rect 20346 12832 20352 12844
rect 20119 12804 20352 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20548 12841 20576 12872
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 17034 12764 17040 12776
rect 16040 12736 17040 12764
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17681 12767 17739 12773
rect 17681 12764 17693 12767
rect 17175 12736 17693 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17681 12733 17693 12736
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 12676 12668 13492 12696
rect 12676 12656 12682 12668
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 16117 12699 16175 12705
rect 16117 12696 16129 12699
rect 13596 12668 16129 12696
rect 13596 12656 13602 12668
rect 16117 12665 16129 12668
rect 16163 12665 16175 12699
rect 16942 12696 16948 12708
rect 16855 12668 16948 12696
rect 16117 12659 16175 12665
rect 16942 12656 16948 12668
rect 17000 12696 17006 12708
rect 17144 12696 17172 12727
rect 17000 12668 17172 12696
rect 17000 12656 17006 12668
rect 9858 12628 9864 12640
rect 9416 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10962 12628 10968 12640
rect 10643 12600 10968 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 12805 12631 12863 12637
rect 12805 12597 12817 12631
rect 12851 12628 12863 12631
rect 13170 12628 13176 12640
rect 12851 12600 13176 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13964 12600 14013 12628
rect 13964 12588 13970 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 14369 12631 14427 12637
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 14458 12628 14464 12640
rect 14415 12600 14464 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 16960 12628 16988 12656
rect 14792 12600 16988 12628
rect 17037 12631 17095 12637
rect 14792 12588 14798 12600
rect 17037 12597 17049 12631
rect 17083 12628 17095 12631
rect 17218 12628 17224 12640
rect 17083 12600 17224 12628
rect 17083 12597 17095 12600
rect 17037 12591 17095 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 18690 12628 18696 12640
rect 18651 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19978 12628 19984 12640
rect 19939 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20622 12628 20628 12640
rect 20583 12600 20628 12628
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 1104 12538 21436 12560
rect 1104 12486 4338 12538
rect 4390 12486 4402 12538
rect 4454 12486 4466 12538
rect 4518 12486 4530 12538
rect 4582 12486 4594 12538
rect 4646 12486 11116 12538
rect 11168 12486 11180 12538
rect 11232 12486 11244 12538
rect 11296 12486 11308 12538
rect 11360 12486 11372 12538
rect 11424 12486 17893 12538
rect 17945 12486 17957 12538
rect 18009 12486 18021 12538
rect 18073 12486 18085 12538
rect 18137 12486 18149 12538
rect 18201 12486 21436 12538
rect 1104 12464 21436 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 1486 12424 1492 12436
rect 1443 12396 1492 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 1486 12384 1492 12396
rect 1544 12384 1550 12436
rect 3142 12424 3148 12436
rect 3103 12396 3148 12424
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 5592 12396 6837 12424
rect 5592 12384 5598 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 6825 12387 6883 12393
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 9490 12424 9496 12436
rect 7340 12396 7788 12424
rect 7340 12384 7346 12396
rect 2869 12359 2927 12365
rect 2869 12325 2881 12359
rect 2915 12356 2927 12359
rect 3786 12356 3792 12368
rect 2915 12328 3792 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 3786 12316 3792 12328
rect 3844 12316 3850 12368
rect 6178 12356 6184 12368
rect 6139 12328 6184 12356
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3050 12288 3056 12300
rect 3007 12260 3056 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 3234 12288 3240 12300
rect 3195 12260 3240 12288
rect 3234 12248 3240 12260
rect 3292 12248 3298 12300
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4948 12260 5089 12288
rect 4948 12248 4954 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5258 12288 5264 12300
rect 5219 12260 5264 12288
rect 5077 12251 5135 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 5408 12260 7021 12288
rect 5408 12248 5414 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7009 12251 7067 12257
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1452 12192 1593 12220
rect 1452 12180 1458 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 1581 12183 1639 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 5994 12220 6000 12232
rect 2823 12192 3004 12220
rect 5955 12192 6000 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 2976 12164 3004 12192
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 6733 12223 6791 12229
rect 6328 12192 6373 12220
rect 6328 12180 6334 12192
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 6822 12220 6828 12232
rect 6779 12192 6828 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7469 12223 7527 12229
rect 7469 12220 7481 12223
rect 7248 12192 7481 12220
rect 7248 12180 7254 12192
rect 7469 12189 7481 12192
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7760 12229 7788 12396
rect 8128 12396 9496 12424
rect 8128 12300 8156 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 11974 12424 11980 12436
rect 11747 12396 11980 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 13446 12424 13452 12436
rect 13407 12396 13452 12424
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 14056 12396 14105 12424
rect 14056 12384 14062 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 15010 12424 15016 12436
rect 14093 12387 14151 12393
rect 14200 12396 15016 12424
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 8260 12328 10241 12356
rect 8260 12316 8266 12328
rect 10229 12325 10241 12328
rect 10275 12356 10287 12359
rect 14200 12356 14228 12396
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15252 12396 15301 12424
rect 15252 12384 15258 12396
rect 15289 12393 15301 12396
rect 15335 12424 15347 12427
rect 16022 12424 16028 12436
rect 15335 12396 16028 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 16022 12384 16028 12396
rect 16080 12384 16086 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 17310 12424 17316 12436
rect 16632 12396 17316 12424
rect 16632 12384 16638 12396
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17678 12424 17684 12436
rect 17635 12396 17684 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 17678 12384 17684 12396
rect 17736 12424 17742 12436
rect 19794 12424 19800 12436
rect 17736 12396 19800 12424
rect 17736 12384 17742 12396
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 19978 12384 19984 12436
rect 20036 12424 20042 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 20036 12396 20085 12424
rect 20036 12384 20042 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 20073 12387 20131 12393
rect 15930 12356 15936 12368
rect 10275 12328 14228 12356
rect 14476 12328 15936 12356
rect 10275 12325 10287 12328
rect 10229 12319 10287 12325
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8110 12288 8116 12300
rect 7975 12260 8116 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 12894 12248 12900 12300
rect 12952 12288 12958 12300
rect 14182 12288 14188 12300
rect 12952 12260 14188 12288
rect 12952 12248 12958 12260
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7616 12192 7665 12220
rect 7616 12180 7622 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12220 10103 12223
rect 10686 12220 10692 12232
rect 10091 12192 10692 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 2958 12112 2964 12164
rect 3016 12112 3022 12164
rect 4985 12155 5043 12161
rect 4985 12121 4997 12155
rect 5031 12152 5043 12155
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5031 12124 5825 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 6288 12152 6316 12180
rect 8036 12152 8064 12183
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10778 12180 10784 12232
rect 10836 12229 10842 12232
rect 10836 12223 10864 12229
rect 10852 12220 10864 12223
rect 11517 12223 11575 12229
rect 10852 12192 11008 12220
rect 10852 12189 10864 12192
rect 10836 12183 10864 12189
rect 10836 12180 10842 12183
rect 6288 12124 8064 12152
rect 10980 12152 11008 12192
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11606 12220 11612 12232
rect 11563 12192 11612 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 12124 12192 12265 12220
rect 12124 12180 12130 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13538 12220 13544 12232
rect 13403 12192 13544 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13964 12192 14105 12220
rect 13964 12180 13970 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 14093 12183 14151 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14476 12220 14504 12328
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 19518 12356 19524 12368
rect 16040 12328 19524 12356
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 15654 12288 15660 12300
rect 14608 12260 15660 12288
rect 14608 12248 14614 12260
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 14415 12192 14504 12220
rect 14645 12223 14703 12229
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 14734 12220 14740 12232
rect 14691 12192 14740 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 13078 12152 13084 12164
rect 10980 12124 13084 12152
rect 5813 12115 5871 12121
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 2133 12087 2191 12093
rect 2133 12053 2145 12087
rect 2179 12084 2191 12087
rect 2590 12084 2596 12096
rect 2179 12056 2596 12084
rect 2179 12053 2191 12056
rect 2133 12047 2191 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 2924 12056 2969 12084
rect 2924 12044 2930 12056
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4120 12056 4629 12084
rect 4120 12044 4126 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4617 12047 4675 12053
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 5408 12056 7021 12084
rect 5408 12044 5414 12056
rect 7009 12053 7021 12056
rect 7055 12053 7067 12087
rect 7009 12047 7067 12053
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 8294 12084 8300 12096
rect 7515 12056 8300 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 10928 12056 10977 12084
rect 10928 12044 10934 12056
rect 10965 12053 10977 12056
rect 11011 12084 11023 12087
rect 14384 12084 14412 12183
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 15105 12223 15163 12229
rect 15105 12220 15117 12223
rect 14884 12192 15117 12220
rect 14884 12180 14890 12192
rect 15105 12189 15117 12192
rect 15151 12189 15163 12223
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15105 12183 15163 12189
rect 15764 12192 15853 12220
rect 15764 12164 15792 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15746 12112 15752 12164
rect 15804 12112 15810 12164
rect 16040 12093 16068 12328
rect 19518 12316 19524 12328
rect 19576 12316 19582 12368
rect 20622 12288 20628 12300
rect 17696 12260 20628 12288
rect 17696 12232 17724 12260
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16264 12192 16681 12220
rect 16264 12180 16270 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16908 12192 17141 12220
rect 16908 12180 16914 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17129 12183 17187 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17678 12220 17684 12232
rect 17460 12192 17505 12220
rect 17591 12192 17684 12220
rect 17460 12180 17466 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 17920 12192 18153 12220
rect 17920 12180 17926 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 19760 12192 20269 12220
rect 19760 12180 19766 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20404 12192 20545 12220
rect 20404 12180 20410 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 19429 12155 19487 12161
rect 19429 12152 19441 12155
rect 16500 12124 19441 12152
rect 16500 12093 16528 12124
rect 19429 12121 19441 12124
rect 19475 12121 19487 12155
rect 19429 12115 19487 12121
rect 19886 12112 19892 12164
rect 19944 12152 19950 12164
rect 20441 12155 20499 12161
rect 20441 12152 20453 12155
rect 19944 12124 20453 12152
rect 19944 12112 19950 12124
rect 20441 12121 20453 12124
rect 20487 12121 20499 12155
rect 20441 12115 20499 12121
rect 11011 12056 14412 12084
rect 16025 12087 16083 12093
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 16025 12053 16037 12087
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12053 16543 12087
rect 16485 12047 16543 12053
rect 17129 12087 17187 12093
rect 17129 12053 17141 12087
rect 17175 12084 17187 12087
rect 17494 12084 17500 12096
rect 17175 12056 17500 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 18196 12056 18245 12084
rect 18196 12044 18202 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 19300 12056 19533 12084
rect 19300 12044 19306 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 1104 11994 21436 12016
rect 1104 11942 7727 11994
rect 7779 11942 7791 11994
rect 7843 11942 7855 11994
rect 7907 11942 7919 11994
rect 7971 11942 7983 11994
rect 8035 11942 14504 11994
rect 14556 11942 14568 11994
rect 14620 11942 14632 11994
rect 14684 11942 14696 11994
rect 14748 11942 14760 11994
rect 14812 11942 21436 11994
rect 1104 11920 21436 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 2188 11852 2329 11880
rect 2188 11840 2194 11852
rect 2317 11849 2329 11852
rect 2363 11880 2375 11883
rect 2682 11880 2688 11892
rect 2363 11852 2688 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 4893 11883 4951 11889
rect 4893 11849 4905 11883
rect 4939 11849 4951 11883
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 4893 11843 4951 11849
rect 3878 11812 3884 11824
rect 3528 11784 3884 11812
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 2314 11747 2372 11753
rect 2314 11713 2326 11747
rect 2360 11744 2372 11747
rect 2682 11744 2688 11756
rect 2360 11716 2544 11744
rect 2643 11716 2688 11744
rect 2360 11713 2372 11716
rect 2314 11707 2372 11713
rect 2516 11676 2544 11716
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 2866 11744 2872 11756
rect 2823 11716 2872 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 2792 11676 2820 11707
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 3528 11753 3556 11784
rect 3878 11772 3884 11784
rect 3936 11812 3942 11824
rect 4908 11812 4936 11843
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 11698 11880 11704 11892
rect 8720 11852 11704 11880
rect 8720 11840 8726 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 12584 11852 14841 11880
rect 12584 11840 12590 11852
rect 14829 11849 14841 11852
rect 14875 11880 14887 11883
rect 15194 11880 15200 11892
rect 14875 11852 15200 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15344 11852 15393 11880
rect 15344 11840 15350 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 16850 11880 16856 11892
rect 16811 11852 16856 11880
rect 15381 11843 15439 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 19150 11880 19156 11892
rect 19107 11852 19156 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 19150 11840 19156 11852
rect 19208 11840 19214 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19576 11852 20484 11880
rect 19576 11840 19582 11852
rect 3936 11784 4936 11812
rect 3936 11772 3942 11784
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 9217 11815 9275 11821
rect 7156 11784 9168 11812
rect 7156 11772 7162 11784
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3970 11744 3976 11756
rect 3835 11716 3976 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 2516 11648 2820 11676
rect 3436 11676 3464 11707
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 4120 11716 4261 11744
rect 4120 11704 4126 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 5307 11716 6377 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6546 11744 6552 11756
rect 6507 11716 6552 11744
rect 6365 11707 6423 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 4798 11676 4804 11688
rect 3436 11648 4804 11676
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 5408 11648 5457 11676
rect 5408 11636 5414 11648
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6236 11648 6745 11676
rect 6236 11636 6242 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 8389 11679 8447 11685
rect 6880 11648 6925 11676
rect 6880 11636 6886 11648
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 8389 11639 8447 11645
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 8404 11608 8432 11639
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 9140 11676 9168 11784
rect 9217 11781 9229 11815
rect 9263 11812 9275 11815
rect 9766 11812 9772 11824
rect 9263 11784 9772 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 9861 11815 9919 11821
rect 9861 11781 9873 11815
rect 9907 11812 9919 11815
rect 10134 11812 10140 11824
rect 9907 11784 10140 11812
rect 9907 11781 9919 11784
rect 9861 11775 9919 11781
rect 10134 11772 10140 11784
rect 10192 11772 10198 11824
rect 15102 11812 15108 11824
rect 12084 11784 13308 11812
rect 12084 11756 12112 11784
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10551 11747 10609 11753
rect 10551 11744 10563 11747
rect 9364 11716 10563 11744
rect 9364 11704 9370 11716
rect 10551 11713 10563 11716
rect 10597 11713 10609 11747
rect 10551 11707 10609 11713
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10410 11676 10416 11688
rect 9140 11648 10416 11676
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 2179 11580 8432 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 9122 11568 9128 11620
rect 9180 11608 9186 11620
rect 10704 11608 10732 11707
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10928 11716 11529 11744
rect 10928 11704 10934 11716
rect 11517 11713 11529 11716
rect 11563 11744 11575 11747
rect 12066 11744 12072 11756
rect 11563 11716 12072 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 12268 11676 12296 11707
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 13280 11753 13308 11784
rect 14016 11784 15108 11812
rect 14016 11753 14044 11784
rect 15102 11772 15108 11784
rect 15160 11772 15166 11824
rect 18138 11772 18144 11824
rect 18196 11812 18202 11824
rect 18966 11812 18972 11824
rect 18196 11784 18972 11812
rect 18196 11772 18202 11784
rect 18966 11772 18972 11784
rect 19024 11812 19030 11824
rect 19024 11784 19656 11812
rect 19024 11772 19030 11784
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12768 11716 13001 11744
rect 12768 11704 12774 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13587 11716 14013 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14642 11744 14648 11756
rect 14555 11716 14648 11744
rect 14001 11707 14059 11713
rect 12894 11676 12900 11688
rect 11020 11648 12900 11676
rect 11020 11636 11026 11648
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 13188 11676 13216 11707
rect 14642 11704 14648 11716
rect 14700 11744 14706 11756
rect 14826 11744 14832 11756
rect 14700 11716 14832 11744
rect 14700 11704 14706 11716
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 15436 11716 15761 11744
rect 15436 11704 15442 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 16298 11744 16304 11756
rect 15749 11707 15807 11713
rect 15948 11716 16304 11744
rect 13188 11648 13308 11676
rect 12250 11608 12256 11620
rect 9180 11580 12256 11608
rect 9180 11568 9186 11580
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 13280 11608 13308 11648
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15344 11648 15853 11676
rect 15344 11636 15350 11648
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 15841 11639 15899 11645
rect 13630 11608 13636 11620
rect 13280 11580 13636 11608
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 15948 11608 15976 11716
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 17405 11747 17463 11753
rect 17405 11744 17417 11747
rect 16356 11716 17417 11744
rect 16356 11704 16362 11716
rect 17405 11713 17417 11716
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17678 11744 17684 11756
rect 17635 11716 17684 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 18233 11747 18291 11753
rect 18233 11744 18245 11747
rect 17828 11716 18245 11744
rect 17828 11704 17834 11716
rect 18233 11713 18245 11716
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 18506 11744 18512 11756
rect 18380 11716 18512 11744
rect 18380 11704 18386 11716
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 18598 11704 18604 11756
rect 18656 11744 18662 11756
rect 19628 11753 19656 11784
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20456 11821 20484 11852
rect 20257 11815 20315 11821
rect 20257 11812 20269 11815
rect 20220 11784 20269 11812
rect 20220 11772 20226 11784
rect 20257 11781 20269 11784
rect 20303 11781 20315 11815
rect 20257 11775 20315 11781
rect 20441 11815 20499 11821
rect 20441 11781 20453 11815
rect 20487 11812 20499 11815
rect 20530 11812 20536 11824
rect 20487 11784 20536 11812
rect 20487 11781 20499 11784
rect 20441 11775 20499 11781
rect 20530 11772 20536 11784
rect 20588 11772 20594 11824
rect 19245 11747 19303 11753
rect 19245 11744 19257 11747
rect 18656 11716 19257 11744
rect 18656 11704 18662 11716
rect 19245 11713 19257 11716
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 18138 11676 18144 11688
rect 17175 11648 18144 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 15304 11580 15976 11608
rect 16040 11608 16068 11639
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 19352 11676 19380 11707
rect 18708 11648 19380 11676
rect 18708 11620 18736 11648
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 20312 11648 20637 11676
rect 20312 11636 20318 11648
rect 20625 11645 20637 11648
rect 20671 11645 20683 11679
rect 20625 11639 20683 11645
rect 16850 11608 16856 11620
rect 16040 11580 16856 11608
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 2924 11512 3249 11540
rect 2924 11500 2930 11512
rect 3237 11509 3249 11512
rect 3283 11509 3295 11543
rect 3237 11503 3295 11509
rect 3697 11543 3755 11549
rect 3697 11509 3709 11543
rect 3743 11540 3755 11543
rect 4154 11540 4160 11552
rect 3743 11512 4160 11540
rect 3743 11509 3755 11512
rect 3697 11503 3755 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4304 11512 4353 11540
rect 4304 11500 4310 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7708 11512 7941 11540
rect 7708 11500 7714 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 8996 11512 9321 11540
rect 8996 11500 9002 11512
rect 9309 11509 9321 11512
rect 9355 11540 9367 11543
rect 9582 11540 9588 11552
rect 9355 11512 9588 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12986 11540 12992 11552
rect 12492 11512 12537 11540
rect 12947 11512 12992 11540
rect 12492 11500 12498 11512
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13136 11512 13461 11540
rect 13136 11500 13142 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 14090 11540 14096 11552
rect 14051 11512 14096 11540
rect 13449 11503 13507 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 15304 11540 15332 11580
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 16908 11580 17325 11608
rect 16908 11568 16914 11580
rect 17313 11577 17325 11580
rect 17359 11577 17371 11611
rect 17313 11571 17371 11577
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 17678 11608 17684 11620
rect 17460 11580 17684 11608
rect 17460 11568 17466 11580
rect 17678 11568 17684 11580
rect 17736 11608 17742 11620
rect 17862 11608 17868 11620
rect 17736 11580 17868 11608
rect 17736 11568 17742 11580
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 18690 11608 18696 11620
rect 18555 11580 18696 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 14608 11512 15332 11540
rect 14608 11500 14614 11512
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 15712 11512 17233 11540
rect 15712 11500 15718 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 17586 11500 17592 11552
rect 17644 11540 17650 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17644 11512 18061 11540
rect 17644 11500 17650 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 19518 11540 19524 11552
rect 19479 11512 19524 11540
rect 18049 11503 18107 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 1104 11450 21436 11472
rect 1104 11398 4338 11450
rect 4390 11398 4402 11450
rect 4454 11398 4466 11450
rect 4518 11398 4530 11450
rect 4582 11398 4594 11450
rect 4646 11398 11116 11450
rect 11168 11398 11180 11450
rect 11232 11398 11244 11450
rect 11296 11398 11308 11450
rect 11360 11398 11372 11450
rect 11424 11398 17893 11450
rect 17945 11398 17957 11450
rect 18009 11398 18021 11450
rect 18073 11398 18085 11450
rect 18137 11398 18149 11450
rect 18201 11398 21436 11450
rect 1104 11376 21436 11398
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11305 2559 11339
rect 2501 11299 2559 11305
rect 2516 11268 2544 11299
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 2740 11308 3801 11336
rect 2740 11296 2746 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 3789 11299 3847 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4706 11296 4712 11348
rect 4764 11296 4770 11348
rect 5997 11339 6055 11345
rect 5997 11305 6009 11339
rect 6043 11336 6055 11339
rect 6270 11336 6276 11348
rect 6043 11308 6276 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 7190 11336 7196 11348
rect 7151 11308 7196 11336
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 9364 11308 9505 11336
rect 9364 11296 9370 11308
rect 9493 11305 9505 11308
rect 9539 11305 9551 11339
rect 10318 11336 10324 11348
rect 9493 11299 9551 11305
rect 9646 11308 10324 11336
rect 3694 11268 3700 11280
rect 2516 11240 3700 11268
rect 3694 11228 3700 11240
rect 3752 11228 3758 11280
rect 4724 11268 4752 11296
rect 6733 11271 6791 11277
rect 6733 11268 6745 11271
rect 4724 11240 6745 11268
rect 6733 11237 6745 11240
rect 6779 11237 6791 11271
rect 6733 11231 6791 11237
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 6972 11240 7665 11268
rect 6972 11228 6978 11240
rect 7653 11237 7665 11240
rect 7699 11237 7711 11271
rect 7653 11231 7711 11237
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 9646 11268 9674 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10962 11336 10968 11348
rect 10744 11308 10968 11336
rect 10744 11296 10750 11308
rect 10962 11296 10968 11308
rect 11020 11336 11026 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 11020 11308 11253 11336
rect 11020 11296 11026 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 12066 11336 12072 11348
rect 11572 11308 12072 11336
rect 11572 11296 11578 11308
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 13044 11308 13093 11336
rect 13044 11296 13050 11308
rect 13081 11305 13093 11308
rect 13127 11336 13139 11339
rect 13446 11336 13452 11348
rect 13127 11308 13452 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14826 11336 14832 11348
rect 14787 11308 14832 11336
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 15528 11308 16589 11336
rect 15528 11296 15534 11308
rect 16577 11305 16589 11308
rect 16623 11336 16635 11339
rect 17770 11336 17776 11348
rect 16623 11308 17776 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 14642 11268 14648 11280
rect 8812 11240 9674 11268
rect 12820 11240 14648 11268
rect 8812 11228 8818 11240
rect 2866 11200 2872 11212
rect 1412 11172 2872 11200
rect 1412 11141 1440 11172
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4706 11200 4712 11212
rect 3988 11172 4292 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1535 11104 2329 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 2317 11101 2329 11104
rect 2363 11132 2375 11135
rect 2406 11132 2412 11144
rect 2363 11104 2412 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 2556 11104 2601 11132
rect 2556 11092 2562 11104
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3988 11141 4016 11172
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 2832 11104 3985 11132
rect 2832 11092 2838 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4120 11104 4213 11132
rect 4120 11092 4126 11104
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 2222 11064 2228 11076
rect 2087 11036 2228 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 2222 11024 2228 11036
rect 2280 11064 2286 11076
rect 2700 11064 2728 11092
rect 2280 11036 2728 11064
rect 2280 11024 2286 11036
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 4080 11064 4108 11092
rect 3384 11036 4108 11064
rect 4264 11064 4292 11172
rect 4356 11172 4712 11200
rect 4356 11141 4384 11172
rect 4706 11160 4712 11172
rect 4764 11200 4770 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4764 11172 4905 11200
rect 4764 11160 4770 11172
rect 4893 11169 4905 11172
rect 4939 11200 4951 11203
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 4939 11172 7481 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 7616 11172 7661 11200
rect 9324 11172 11284 11200
rect 7616 11160 7622 11172
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5626 11132 5632 11144
rect 4847 11104 5632 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 4816 11064 4844 11095
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5868 11104 5917 11132
rect 5868 11092 5874 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 5905 11095 5963 11101
rect 6012 11104 6561 11132
rect 4264 11036 4844 11064
rect 3384 11024 3390 11036
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 6012 11064 6040 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 7190 11092 7196 11144
rect 7248 11132 7254 11144
rect 7650 11132 7656 11144
rect 7248 11104 7656 11132
rect 7248 11092 7254 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 5776 11036 6040 11064
rect 5776 11024 5782 11036
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 7944 11064 7972 11095
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9324 11141 9352 11172
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9180 11104 9321 11132
rect 9180 11092 9186 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9824 11104 10149 11132
rect 9824 11092 9830 11104
rect 10137 11101 10149 11104
rect 10183 11132 10195 11135
rect 10778 11132 10784 11144
rect 10183 11104 10784 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11256 11141 11284 11172
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 12342 11132 12348 11144
rect 11471 11104 12348 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 12342 11092 12348 11104
rect 12400 11132 12406 11144
rect 12820 11132 12848 11240
rect 14642 11228 14648 11240
rect 14700 11228 14706 11280
rect 16022 11268 16028 11280
rect 15580 11240 16028 11268
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13173 11203 13231 11209
rect 12952 11172 13124 11200
rect 12952 11160 12958 11172
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12400 11104 13001 11132
rect 12400 11092 12406 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 13096 11132 13124 11172
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 14090 11200 14096 11212
rect 13219 11172 14096 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 14090 11160 14096 11172
rect 14148 11200 14154 11212
rect 14921 11203 14979 11209
rect 14148 11172 14872 11200
rect 14148 11160 14154 11172
rect 13262 11132 13268 11144
rect 13096 11104 13268 11132
rect 12989 11095 13047 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13630 11132 13636 11144
rect 13495 11104 13636 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 14660 11141 14688 11172
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14844 11132 14872 11172
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 15286 11200 15292 11212
rect 14967 11172 15292 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15580 11209 15608 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 16908 11240 17724 11268
rect 16908 11228 16914 11240
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 15838 11200 15844 11212
rect 15703 11172 15844 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 17586 11200 17592 11212
rect 15948 11172 16712 11200
rect 17547 11172 17592 11200
rect 15948 11132 15976 11172
rect 14844 11104 15976 11132
rect 16032 11135 16090 11141
rect 14737 11095 14795 11101
rect 16032 11101 16044 11135
rect 16078 11132 16090 11135
rect 16298 11132 16304 11144
rect 16078 11104 16304 11132
rect 16078 11101 16090 11104
rect 16032 11095 16090 11101
rect 6328 11036 7972 11064
rect 6328 11024 6334 11036
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 9582 11064 9588 11076
rect 8628 11036 9588 11064
rect 8628 11024 8634 11036
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 14550 11064 14556 11076
rect 12492 11036 14556 11064
rect 12492 11024 12498 11036
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14752 11064 14780 11095
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 16684 11141 16712 11172
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 17696 11209 17724 11240
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11200 17739 11203
rect 17727 11172 19104 11200
rect 17727 11169 17739 11172
rect 17681 11163 17739 11169
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 14826 11064 14832 11076
rect 14739 11036 14832 11064
rect 14826 11024 14832 11036
rect 14884 11064 14890 11076
rect 16500 11064 16528 11095
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17126 11132 17132 11144
rect 16816 11104 17132 11132
rect 16816 11092 16822 11104
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17494 11132 17500 11144
rect 17455 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18509 11135 18567 11141
rect 18509 11101 18521 11135
rect 18555 11132 18567 11135
rect 18966 11132 18972 11144
rect 18555 11104 18972 11132
rect 18555 11101 18567 11104
rect 18509 11095 18567 11101
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 19076 11132 19104 11172
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19794 11200 19800 11212
rect 19392 11172 19800 11200
rect 19392 11160 19398 11172
rect 19794 11160 19800 11172
rect 19852 11200 19858 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19852 11172 20177 11200
rect 19852 11160 19858 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 19426 11132 19432 11144
rect 19076 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 17586 11064 17592 11076
rect 14884 11036 16528 11064
rect 17144 11036 17592 11064
rect 14884 11024 14890 11036
rect 2682 10996 2688 11008
rect 2643 10968 2688 10996
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 6972 10968 7849 10996
rect 6972 10956 6978 10968
rect 7837 10965 7849 10968
rect 7883 10996 7895 10999
rect 8202 10996 8208 11008
rect 7883 10968 8208 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 11606 10996 11612 11008
rect 11519 10968 11612 10996
rect 11606 10956 11612 10968
rect 11664 10996 11670 11008
rect 12250 10996 12256 11008
rect 11664 10968 12256 10996
rect 11664 10956 11670 10968
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 15654 10996 15660 11008
rect 15252 10968 15660 10996
rect 15252 10956 15258 10968
rect 15654 10956 15660 10968
rect 15712 10996 15718 11008
rect 15749 10999 15807 11005
rect 15749 10996 15761 10999
rect 15712 10968 15761 10996
rect 15712 10956 15718 10968
rect 15749 10965 15761 10968
rect 15795 10965 15807 10999
rect 15749 10959 15807 10965
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 16390 10996 16396 11008
rect 15988 10968 16396 10996
rect 15988 10956 15994 10968
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17144 11005 17172 11036
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 18690 11064 18696 11076
rect 18651 11036 18696 11064
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 17129 10999 17187 11005
rect 17129 10965 17141 10999
rect 17175 10965 17187 10999
rect 17129 10959 17187 10965
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19613 10999 19671 11005
rect 19613 10996 19625 10999
rect 19392 10968 19625 10996
rect 19392 10956 19398 10968
rect 19613 10965 19625 10968
rect 19659 10965 19671 10999
rect 19978 10996 19984 11008
rect 19939 10968 19984 10996
rect 19613 10959 19671 10965
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 20070 10956 20076 11008
rect 20128 10996 20134 11008
rect 20128 10968 20173 10996
rect 20128 10956 20134 10968
rect 1104 10906 21436 10928
rect 1104 10854 7727 10906
rect 7779 10854 7791 10906
rect 7843 10854 7855 10906
rect 7907 10854 7919 10906
rect 7971 10854 7983 10906
rect 8035 10854 14504 10906
rect 14556 10854 14568 10906
rect 14620 10854 14632 10906
rect 14684 10854 14696 10906
rect 14748 10854 14760 10906
rect 14812 10854 21436 10906
rect 1104 10832 21436 10854
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 2498 10792 2504 10804
rect 2096 10764 2504 10792
rect 2096 10752 2102 10764
rect 2498 10752 2504 10764
rect 2556 10792 2562 10804
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2556 10764 2697 10792
rect 2556 10752 2562 10764
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 3970 10792 3976 10804
rect 2685 10755 2743 10761
rect 3528 10764 3976 10792
rect 2222 10684 2228 10736
rect 2280 10724 2286 10736
rect 2317 10727 2375 10733
rect 2317 10724 2329 10727
rect 2280 10696 2329 10724
rect 2280 10684 2286 10696
rect 2317 10693 2329 10696
rect 2363 10693 2375 10727
rect 2317 10687 2375 10693
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10724 2467 10727
rect 2774 10724 2780 10736
rect 2455 10696 2780 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3528 10724 3556 10764
rect 3970 10752 3976 10764
rect 4028 10792 4034 10804
rect 4028 10764 4568 10792
rect 4028 10752 4034 10764
rect 4249 10727 4307 10733
rect 4249 10724 4261 10727
rect 3436 10696 3556 10724
rect 3620 10696 4261 10724
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 1489 10619 1547 10625
rect 1504 10520 1532 10619
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 3326 10656 3332 10668
rect 2547 10628 3332 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 3436 10665 3464 10696
rect 3620 10665 3648 10696
rect 4249 10693 4261 10696
rect 4295 10693 4307 10727
rect 4249 10687 4307 10693
rect 4540 10724 4568 10764
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5626 10792 5632 10804
rect 4856 10764 5632 10792
rect 4856 10752 4862 10764
rect 5626 10752 5632 10764
rect 5684 10792 5690 10804
rect 7650 10792 7656 10804
rect 5684 10764 7656 10792
rect 5684 10752 5690 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8720 10764 9505 10792
rect 8720 10752 8726 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 14737 10795 14795 10801
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 14826 10792 14832 10804
rect 14783 10764 14832 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15841 10795 15899 10801
rect 15841 10761 15853 10795
rect 15887 10792 15899 10795
rect 16298 10792 16304 10804
rect 15887 10764 16304 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 19978 10792 19984 10804
rect 19659 10764 19984 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 6365 10727 6423 10733
rect 4540 10696 5764 10724
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 3526 10659 3584 10665
rect 3526 10625 3538 10659
rect 3572 10625 3584 10659
rect 3620 10659 3684 10665
rect 3620 10628 3638 10659
rect 3526 10619 3584 10625
rect 3626 10625 3638 10628
rect 3672 10625 3684 10659
rect 3786 10656 3792 10668
rect 3747 10628 3792 10656
rect 3626 10619 3684 10625
rect 3528 10588 3556 10619
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4540 10665 4568 10696
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4212 10628 4445 10656
rect 4212 10616 4218 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4525 10619 4583 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 5626 10656 5632 10668
rect 5587 10628 5632 10656
rect 4801 10619 4859 10625
rect 4172 10588 4200 10616
rect 3528 10560 4200 10588
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4816 10588 4844 10619
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 5736 10665 5764 10696
rect 6365 10693 6377 10727
rect 6411 10724 6423 10727
rect 8938 10724 8944 10736
rect 6411 10696 7604 10724
rect 6411 10693 6423 10696
rect 6365 10687 6423 10693
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 5767 10628 6653 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6641 10619 6699 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7576 10665 7604 10696
rect 7852 10696 8944 10724
rect 7852 10668 7880 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 12802 10724 12808 10736
rect 12763 10696 12808 10724
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 13538 10684 13544 10736
rect 13596 10724 13602 10736
rect 15473 10727 15531 10733
rect 13596 10696 14504 10724
rect 13596 10684 13602 10696
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 4304 10560 4844 10588
rect 4304 10548 4310 10560
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7116 10588 7144 10619
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7708 10628 7757 10656
rect 7708 10616 7714 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8113 10659 8171 10665
rect 7892 10628 7937 10656
rect 7892 10616 7898 10628
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 8128 10588 8156 10619
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8260 10628 8585 10656
rect 8260 10616 8266 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 10042 10656 10048 10668
rect 10003 10628 10048 10656
rect 9309 10619 9367 10625
rect 6880 10560 8156 10588
rect 6880 10548 6886 10560
rect 9214 10548 9220 10600
rect 9272 10548 9278 10600
rect 9324 10588 9352 10619
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10744 10628 10793 10656
rect 10744 10616 10750 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12986 10656 12992 10668
rect 12023 10628 12992 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14476 10665 14504 10696
rect 15473 10693 15485 10727
rect 15519 10724 15531 10727
rect 16114 10724 16120 10736
rect 15519 10696 16120 10724
rect 15519 10693 15531 10696
rect 15473 10687 15531 10693
rect 16114 10684 16120 10696
rect 16172 10684 16178 10736
rect 17957 10727 18015 10733
rect 17957 10693 17969 10727
rect 18003 10724 18015 10727
rect 18598 10724 18604 10736
rect 18003 10696 18604 10724
rect 18003 10693 18015 10696
rect 17957 10687 18015 10693
rect 18598 10684 18604 10696
rect 18656 10684 18662 10736
rect 19334 10724 19340 10736
rect 18800 10696 19340 10724
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14642 10656 14648 10668
rect 14507 10628 14648 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 16666 10656 16672 10668
rect 16627 10628 16672 10656
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 18800 10665 18828 10696
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17828 10628 17877 10656
rect 17828 10616 17834 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 19058 10656 19064 10668
rect 19019 10628 19064 10656
rect 18785 10619 18843 10625
rect 10870 10588 10876 10600
rect 9324 10560 10876 10588
rect 10870 10548 10876 10560
rect 10928 10588 10934 10600
rect 11698 10588 11704 10600
rect 10928 10560 11704 10588
rect 10928 10548 10934 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 13630 10548 13636 10600
rect 13688 10588 13694 10600
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 13688 10560 14749 10588
rect 13688 10548 13694 10560
rect 14737 10557 14749 10560
rect 14783 10557 14795 10591
rect 14737 10551 14795 10557
rect 8938 10520 8944 10532
rect 1504 10492 8944 10520
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 9232 10520 9260 10548
rect 9858 10520 9864 10532
rect 9232 10492 9864 10520
rect 9858 10480 9864 10492
rect 9916 10520 9922 10532
rect 10229 10523 10287 10529
rect 10229 10520 10241 10523
rect 9916 10492 10241 10520
rect 9916 10480 9922 10492
rect 10229 10489 10241 10492
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 13722 10520 13728 10532
rect 10468 10492 13728 10520
rect 10468 10480 10474 10492
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 14001 10523 14059 10529
rect 14001 10489 14013 10523
rect 14047 10520 14059 10523
rect 14182 10520 14188 10532
rect 14047 10492 14188 10520
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 14752 10520 14780 10551
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18708 10588 18736 10619
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19668 10628 19809 10656
rect 19668 10616 19674 10628
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 20530 10656 20536 10668
rect 20491 10628 20536 10656
rect 19797 10619 19855 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 17736 10560 18736 10588
rect 18969 10591 19027 10597
rect 17736 10548 17742 10560
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19518 10588 19524 10600
rect 19015 10560 19524 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 20036 10560 20085 10588
rect 20036 10548 20042 10560
rect 20073 10557 20085 10560
rect 20119 10588 20131 10591
rect 20622 10588 20628 10600
rect 20119 10560 20628 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 14752 10492 20668 10520
rect 20640 10464 20668 10492
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3016 10424 3157 10452
rect 3016 10412 3022 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 6733 10455 6791 10461
rect 6733 10452 6745 10455
rect 6696 10424 6745 10452
rect 6696 10412 6702 10424
rect 6733 10421 6745 10424
rect 6779 10421 6791 10455
rect 6733 10415 6791 10421
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 7558 10452 7564 10464
rect 6880 10424 6925 10452
rect 7519 10424 7564 10452
rect 6880 10412 6886 10424
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7708 10424 8033 10452
rect 7708 10412 7714 10424
rect 8021 10421 8033 10424
rect 8067 10452 8079 10455
rect 8110 10452 8116 10464
rect 8067 10424 8116 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 8110 10412 8116 10424
rect 8168 10452 8174 10464
rect 8662 10452 8668 10464
rect 8168 10424 8668 10452
rect 8168 10412 8174 10424
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8757 10455 8815 10461
rect 8757 10421 8769 10455
rect 8803 10452 8815 10455
rect 9214 10452 9220 10464
rect 8803 10424 9220 10452
rect 8803 10421 8815 10424
rect 8757 10415 8815 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10652 10424 10885 10452
rect 10652 10412 10658 10424
rect 10873 10421 10885 10424
rect 10919 10421 10931 10455
rect 14550 10452 14556 10464
rect 14511 10424 14556 10452
rect 10873 10415 10931 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 16482 10452 16488 10464
rect 15896 10424 16488 10452
rect 15896 10412 15902 10424
rect 16482 10412 16488 10424
rect 16540 10452 16546 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16540 10424 16773 10452
rect 16540 10412 16546 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 19610 10452 19616 10464
rect 17276 10424 19616 10452
rect 17276 10412 17282 10424
rect 19610 10412 19616 10424
rect 19668 10412 19674 10464
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 19981 10455 20039 10461
rect 19981 10452 19993 10455
rect 19944 10424 19993 10452
rect 19944 10412 19950 10424
rect 19981 10421 19993 10424
rect 20027 10421 20039 10455
rect 20622 10452 20628 10464
rect 20583 10424 20628 10452
rect 19981 10415 20039 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 1104 10362 21436 10384
rect 1104 10310 4338 10362
rect 4390 10310 4402 10362
rect 4454 10310 4466 10362
rect 4518 10310 4530 10362
rect 4582 10310 4594 10362
rect 4646 10310 11116 10362
rect 11168 10310 11180 10362
rect 11232 10310 11244 10362
rect 11296 10310 11308 10362
rect 11360 10310 11372 10362
rect 11424 10310 17893 10362
rect 17945 10310 17957 10362
rect 18009 10310 18021 10362
rect 18073 10310 18085 10362
rect 18137 10310 18149 10362
rect 18201 10310 21436 10362
rect 1104 10288 21436 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2556 10220 2789 10248
rect 2556 10208 2562 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4154 10248 4160 10260
rect 4019 10220 4160 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7834 10248 7840 10260
rect 7340 10220 7840 10248
rect 7340 10208 7346 10220
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8938 10248 8944 10260
rect 8352 10220 8397 10248
rect 8899 10220 8944 10248
rect 8352 10208 8358 10220
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9398 10248 9404 10260
rect 9324 10220 9404 10248
rect 4709 10183 4767 10189
rect 4709 10149 4721 10183
rect 4755 10180 4767 10183
rect 6454 10180 6460 10192
rect 4755 10152 6460 10180
rect 4755 10149 4767 10152
rect 4709 10143 4767 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6972 10084 7021 10112
rect 6972 10072 6978 10084
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 9324 10112 9352 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 10042 10248 10048 10260
rect 9548 10220 10048 10248
rect 9548 10208 9554 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10468 10220 10609 10248
rect 10468 10208 10474 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 12342 10248 12348 10260
rect 10735 10220 12348 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12618 10248 12624 10260
rect 12483 10220 12624 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13262 10248 13268 10260
rect 13219 10220 13268 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 13780 10220 14504 10248
rect 13780 10208 13786 10220
rect 10781 10183 10839 10189
rect 10781 10149 10793 10183
rect 10827 10180 10839 10183
rect 12986 10180 12992 10192
rect 10827 10152 12992 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 14476 10180 14504 10220
rect 14550 10208 14556 10260
rect 14608 10248 14614 10260
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 14608 10220 16129 10248
rect 14608 10208 14614 10220
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 19337 10251 19395 10257
rect 16117 10211 16175 10217
rect 16408 10220 18092 10248
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 14476 10152 15485 10180
rect 15473 10149 15485 10152
rect 15519 10180 15531 10183
rect 16408 10180 16436 10220
rect 15519 10152 16436 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 16482 10140 16488 10192
rect 16540 10180 16546 10192
rect 18064 10180 18092 10220
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19518 10248 19524 10260
rect 19383 10220 19524 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 19886 10248 19892 10260
rect 19625 10220 19892 10248
rect 19625 10180 19653 10220
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20070 10248 20076 10260
rect 20031 10220 20076 10248
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 19978 10180 19984 10192
rect 16540 10152 17448 10180
rect 18064 10152 19653 10180
rect 19939 10152 19984 10180
rect 16540 10140 16546 10152
rect 9401 10115 9459 10121
rect 9401 10112 9413 10115
rect 9324 10084 9413 10112
rect 7009 10075 7067 10081
rect 9401 10081 9413 10084
rect 9447 10081 9459 10115
rect 9582 10112 9588 10124
rect 9543 10084 9588 10112
rect 9401 10075 9459 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16724 10084 17356 10112
rect 16724 10072 16730 10084
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 2464 10016 2513 10044
rect 2464 10004 2470 10016
rect 2501 10013 2513 10016
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 2866 10044 2872 10056
rect 2648 10016 2693 10044
rect 2827 10016 2872 10044
rect 2648 10004 2654 10016
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3878 10044 3884 10056
rect 3839 10016 3884 10044
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 5074 10044 5080 10056
rect 4571 10016 5080 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5442 10044 5448 10056
rect 5399 10016 5448 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5626 10044 5632 10056
rect 5583 10016 5632 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7558 10044 7564 10056
rect 6871 10016 7564 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 8168 10016 8217 10044
rect 8168 10004 8174 10016
rect 8205 10013 8217 10016
rect 8251 10013 8263 10047
rect 10870 10044 10876 10056
rect 10831 10016 10876 10044
rect 8205 10007 8263 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 1670 9976 1676 9988
rect 1631 9948 1676 9976
rect 1670 9936 1676 9948
rect 1728 9936 1734 9988
rect 2317 9979 2375 9985
rect 2317 9945 2329 9979
rect 2363 9976 2375 9979
rect 6917 9979 6975 9985
rect 6917 9976 6929 9979
rect 2363 9948 6929 9976
rect 2363 9945 2375 9948
rect 2317 9939 2375 9945
rect 6917 9945 6929 9948
rect 6963 9945 6975 9979
rect 11072 9976 11100 10007
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11480 10016 11529 10044
rect 11480 10004 11486 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10044 12311 10047
rect 12526 10044 12532 10056
rect 12299 10016 12532 10044
rect 12299 10013 12311 10016
rect 12253 10007 12311 10013
rect 12526 10004 12532 10016
rect 12584 10044 12590 10056
rect 12986 10044 12992 10056
rect 12584 10016 12992 10044
rect 12584 10004 12590 10016
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 11606 9976 11612 9988
rect 6917 9939 6975 9945
rect 10060 9948 11008 9976
rect 11072 9948 11612 9976
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 5442 9908 5448 9920
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6328 9880 6469 9908
rect 6328 9868 6334 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 8996 9880 9321 9908
rect 8996 9868 9002 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10060 9908 10088 9948
rect 9548 9880 10088 9908
rect 9548 9868 9554 9880
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10192 9880 10333 9908
rect 10192 9868 10198 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 10980 9908 11008 9948
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 13188 9976 13216 10007
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 17328 10053 17356 10084
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 13872 10016 15301 10044
rect 13872 10004 13878 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 16025 10047 16083 10053
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17420 10044 17448 10152
rect 19978 10140 19984 10152
rect 20036 10140 20042 10192
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 20165 10115 20223 10121
rect 20165 10081 20177 10115
rect 20211 10112 20223 10115
rect 20254 10112 20260 10124
rect 20211 10084 20260 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 17420 10016 17969 10044
rect 17313 10007 17371 10013
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 14366 9976 14372 9988
rect 13188 9948 14372 9976
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 14642 9976 14648 9988
rect 14603 9948 14648 9976
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 15010 9976 15016 9988
rect 14875 9948 15016 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 15010 9936 15016 9948
rect 15068 9936 15074 9988
rect 16040 9976 16068 10007
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18104 10016 18149 10044
rect 18104 10004 18110 10016
rect 15120 9948 16068 9976
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 10980 9880 11713 9908
rect 10321 9871 10379 9877
rect 11701 9877 11713 9880
rect 11747 9908 11759 9911
rect 13078 9908 13084 9920
rect 11747 9880 13084 9908
rect 11747 9877 11759 9880
rect 11701 9871 11759 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 13722 9908 13728 9920
rect 13403 9880 13728 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 15120 9908 15148 9948
rect 16206 9936 16212 9988
rect 16264 9976 16270 9988
rect 16666 9976 16672 9988
rect 16264 9948 16672 9976
rect 16264 9936 16270 9948
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 17129 9979 17187 9985
rect 17129 9945 17141 9979
rect 17175 9976 17187 9979
rect 17218 9976 17224 9988
rect 17175 9948 17224 9976
rect 17175 9945 17187 9948
rect 17129 9939 17187 9945
rect 17218 9936 17224 9948
rect 17276 9936 17282 9988
rect 17494 9976 17500 9988
rect 17407 9948 17500 9976
rect 17494 9936 17500 9948
rect 17552 9976 17558 9988
rect 18248 9976 18276 10075
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20622 10044 20628 10056
rect 19935 10016 20628 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 17552 9948 18276 9976
rect 17552 9936 17558 9948
rect 18230 9908 18236 9920
rect 14056 9880 15148 9908
rect 18191 9880 18236 9908
rect 14056 9868 14062 9880
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 1104 9818 21436 9840
rect 1104 9766 7727 9818
rect 7779 9766 7791 9818
rect 7843 9766 7855 9818
rect 7907 9766 7919 9818
rect 7971 9766 7983 9818
rect 8035 9766 14504 9818
rect 14556 9766 14568 9818
rect 14620 9766 14632 9818
rect 14684 9766 14696 9818
rect 14748 9766 14760 9818
rect 14812 9766 21436 9818
rect 1104 9744 21436 9766
rect 5442 9704 5448 9716
rect 4724 9676 5448 9704
rect 2958 9636 2964 9648
rect 2332 9608 2964 9636
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 2332 9577 2360 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 4724 9645 4752 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6822 9704 6828 9716
rect 6420 9676 6828 9704
rect 6420 9664 6426 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 8294 9704 8300 9716
rect 6972 9676 8300 9704
rect 6972 9664 6978 9676
rect 4709 9639 4767 9645
rect 4709 9605 4721 9639
rect 4755 9605 4767 9639
rect 4709 9599 4767 9605
rect 4893 9639 4951 9645
rect 4893 9605 4905 9639
rect 4939 9636 4951 9639
rect 4939 9608 5672 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 5644 9580 5672 9608
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7944 9636 7972 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 9548 9676 9781 9704
rect 9548 9664 9554 9676
rect 9769 9673 9781 9676
rect 9815 9673 9827 9707
rect 9769 9667 9827 9673
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 12437 9707 12495 9713
rect 12437 9704 12449 9707
rect 10100 9676 12449 9704
rect 10100 9664 10106 9676
rect 12437 9673 12449 9676
rect 12483 9673 12495 9707
rect 12437 9667 12495 9673
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 13909 9707 13967 9713
rect 13909 9704 13921 9707
rect 13872 9676 13921 9704
rect 13872 9664 13878 9676
rect 13909 9673 13921 9676
rect 13955 9673 13967 9707
rect 13909 9667 13967 9673
rect 14274 9664 14280 9716
rect 14332 9704 14338 9716
rect 17494 9704 17500 9716
rect 14332 9676 17500 9704
rect 14332 9664 14338 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 8570 9636 8576 9648
rect 7156 9608 7604 9636
rect 7944 9608 8576 9636
rect 7156 9596 7162 9608
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1452 9540 1685 9568
rect 1452 9528 1458 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2682 9568 2688 9580
rect 2547 9540 2688 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 1688 9500 1716 9531
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3050 9568 3056 9580
rect 3011 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9568 3114 9580
rect 3418 9568 3424 9580
rect 3108 9540 3424 9568
rect 3108 9528 3114 9540
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5350 9568 5356 9580
rect 5031 9540 5356 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 1762 9500 1768 9512
rect 1688 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 1912 9472 2605 9500
rect 1912 9460 1918 9472
rect 2593 9469 2605 9472
rect 2639 9500 2651 9503
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2639 9472 3157 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 1486 9432 1492 9444
rect 1447 9404 1492 9432
rect 1486 9392 1492 9404
rect 1544 9392 1550 9444
rect 1780 9432 1808 9460
rect 3896 9432 3924 9531
rect 5350 9528 5356 9540
rect 5408 9568 5414 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5408 9540 5457 9568
rect 5408 9528 5414 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 6086 9568 6092 9580
rect 5684 9540 6092 9568
rect 5684 9528 5690 9540
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 7006 9568 7012 9580
rect 6411 9540 7012 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 6380 9500 6408 9531
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7466 9568 7472 9580
rect 7427 9540 7472 9568
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7576 9577 7604 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 12400 9608 14320 9636
rect 12400 9596 12406 9608
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 8720 9540 9522 9568
rect 8720 9528 8726 9540
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11480 9540 11529 9568
rect 11480 9528 11486 9540
rect 11517 9537 11529 9540
rect 11563 9568 11575 9571
rect 12250 9568 12256 9580
rect 11563 9540 12256 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 13538 9568 13544 9580
rect 13499 9540 13544 9568
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 13998 9568 14004 9580
rect 13648 9540 14004 9568
rect 13648 9512 13676 9540
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 14292 9568 14320 9608
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 14424 9608 14473 9636
rect 14424 9596 14430 9608
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17402 9636 17408 9648
rect 17175 9608 17408 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17402 9596 17408 9608
rect 17460 9636 17466 9648
rect 18325 9639 18383 9645
rect 17460 9608 18276 9636
rect 17460 9596 17466 9608
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 14292 9540 14657 9568
rect 14645 9537 14657 9540
rect 14691 9568 14703 9571
rect 15102 9568 15108 9580
rect 14691 9540 15108 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17494 9568 17500 9580
rect 17359 9540 17500 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 5644 9472 6408 9500
rect 5644 9432 5672 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7432 9472 7757 9500
rect 7432 9460 7438 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9030 9500 9036 9512
rect 8803 9472 9036 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 11974 9500 11980 9512
rect 10534 9486 11980 9500
rect 10520 9472 11980 9486
rect 1780 9404 3924 9432
rect 5552 9404 5672 9432
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 4982 9364 4988 9376
rect 4755 9336 4988 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5552 9373 5580 9404
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 7653 9435 7711 9441
rect 7653 9432 7665 9435
rect 6052 9404 7665 9432
rect 6052 9392 6058 9404
rect 7653 9401 7665 9404
rect 7699 9401 7711 9435
rect 7653 9395 7711 9401
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 9582 9432 9588 9444
rect 8352 9404 9588 9432
rect 8352 9392 8358 9404
rect 9582 9392 9588 9404
rect 9640 9432 9646 9444
rect 10520 9432 10548 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 12483 9472 12633 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12621 9469 12633 9472
rect 12667 9500 12679 9503
rect 13630 9500 13636 9512
rect 12667 9472 13636 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 15856 9500 15884 9531
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 18104 9540 18153 9568
rect 18104 9528 18110 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18248 9568 18276 9608
rect 18325 9605 18337 9639
rect 18371 9636 18383 9639
rect 18598 9636 18604 9648
rect 18371 9608 18604 9636
rect 18371 9605 18383 9608
rect 18325 9599 18383 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 18690 9596 18696 9648
rect 18748 9636 18754 9648
rect 18748 9608 19932 9636
rect 18748 9596 18754 9608
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 18248 9540 18429 9568
rect 18141 9531 18199 9537
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 13780 9472 15884 9500
rect 18156 9500 18184 9531
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 19904 9577 19932 9608
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18564 9540 18889 9568
rect 18564 9528 18570 9540
rect 18877 9537 18889 9540
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 19935 9540 20545 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20533 9537 20545 9540
rect 20579 9537 20591 9571
rect 20533 9531 20591 9537
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18156 9472 18981 9500
rect 13780 9460 13786 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19300 9472 20392 9500
rect 19300 9460 19306 9472
rect 9640 9404 10548 9432
rect 11701 9435 11759 9441
rect 9640 9392 9646 9404
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 11790 9432 11796 9444
rect 11747 9404 11796 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 11790 9392 11796 9404
rect 11848 9392 11854 9444
rect 12544 9404 13584 9432
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5813 9367 5871 9373
rect 5813 9364 5825 9367
rect 5684 9336 5825 9364
rect 5684 9324 5690 9336
rect 5813 9333 5825 9336
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6236 9336 6469 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 10410 9364 10416 9376
rect 6880 9336 10416 9364
rect 6880 9324 6886 9336
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10594 9324 10600 9376
rect 10652 9364 10658 9376
rect 12544 9373 12572 9404
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 10652 9336 12541 9364
rect 10652 9324 10658 9336
rect 12529 9333 12541 9336
rect 12575 9364 12587 9367
rect 12618 9364 12624 9376
rect 12575 9336 12624 9364
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13556 9373 13584 9404
rect 17218 9392 17224 9444
rect 17276 9392 17282 9444
rect 17957 9435 18015 9441
rect 17957 9401 17969 9435
rect 18003 9432 18015 9435
rect 19794 9432 19800 9444
rect 18003 9404 19800 9432
rect 18003 9401 18015 9404
rect 17957 9395 18015 9401
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 20364 9441 20392 9472
rect 20349 9435 20407 9441
rect 20349 9401 20361 9435
rect 20395 9401 20407 9435
rect 20349 9395 20407 9401
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12768 9336 12909 9364
rect 12768 9324 12774 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9333 13599 9367
rect 13541 9327 13599 9333
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14884 9336 15301 9364
rect 14884 9324 14890 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16298 9364 16304 9376
rect 16071 9336 16304 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17236 9364 17264 9392
rect 17494 9364 17500 9376
rect 17236 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 19702 9364 19708 9376
rect 19663 9336 19708 9364
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 1104 9274 21436 9296
rect 1104 9222 4338 9274
rect 4390 9222 4402 9274
rect 4454 9222 4466 9274
rect 4518 9222 4530 9274
rect 4582 9222 4594 9274
rect 4646 9222 11116 9274
rect 11168 9222 11180 9274
rect 11232 9222 11244 9274
rect 11296 9222 11308 9274
rect 11360 9222 11372 9274
rect 11424 9222 17893 9274
rect 17945 9222 17957 9274
rect 18009 9222 18021 9274
rect 18073 9222 18085 9274
rect 18137 9222 18149 9274
rect 18201 9222 21436 9274
rect 1104 9200 21436 9222
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 8938 9160 8944 9172
rect 6144 9132 8944 9160
rect 6144 9120 6150 9132
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9548 9132 9965 9160
rect 9548 9120 9554 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 9953 9123 10011 9129
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 14366 9160 14372 9172
rect 10928 9132 14372 9160
rect 10928 9120 10934 9132
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15565 9163 15623 9169
rect 15565 9160 15577 9163
rect 15160 9132 15577 9160
rect 15160 9120 15166 9132
rect 15565 9129 15577 9132
rect 15611 9129 15623 9163
rect 15565 9123 15623 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18506 9160 18512 9172
rect 17552 9132 18512 9160
rect 17552 9120 17558 9132
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 7374 9092 7380 9104
rect 7335 9064 7380 9092
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 12345 9095 12403 9101
rect 12345 9092 12357 9095
rect 10468 9064 12357 9092
rect 10468 9052 10474 9064
rect 12345 9061 12357 9064
rect 12391 9092 12403 9095
rect 15378 9092 15384 9104
rect 12391 9064 15384 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 15378 9052 15384 9064
rect 15436 9092 15442 9104
rect 15657 9095 15715 9101
rect 15657 9092 15669 9095
rect 15436 9064 15669 9092
rect 15436 9052 15442 9064
rect 15657 9061 15669 9064
rect 15703 9061 15715 9095
rect 15657 9055 15715 9061
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 18690 9092 18696 9104
rect 16724 9064 18696 9092
rect 16724 9052 16730 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 3694 9024 3700 9036
rect 1872 8996 3700 9024
rect 1872 8965 1900 8996
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5166 9024 5172 9036
rect 5127 8996 5172 9024
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 6178 9024 6184 9036
rect 5316 8996 6184 9024
rect 5316 8984 5322 8996
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7156 8996 7481 9024
rect 7156 8984 7162 8996
rect 7469 8993 7481 8996
rect 7515 9024 7527 9027
rect 7650 9024 7656 9036
rect 7515 8996 7656 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 10686 9024 10692 9036
rect 8036 8996 10692 9024
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 1857 8919 1915 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3200 8928 3801 8956
rect 3200 8916 3206 8928
rect 3789 8925 3801 8928
rect 3835 8956 3847 8959
rect 4154 8956 4160 8968
rect 3835 8928 4160 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 5902 8956 5908 8968
rect 5863 8928 5908 8956
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6788 8928 7021 8956
rect 6788 8916 6794 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7009 8919 7067 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7561 8959 7619 8965
rect 7340 8928 7433 8956
rect 7340 8916 7346 8928
rect 7561 8925 7573 8959
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 5994 8888 6000 8900
rect 4939 8860 6000 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 7300 8888 7328 8916
rect 6972 8860 7328 8888
rect 6972 8848 6978 8860
rect 7466 8848 7472 8900
rect 7524 8888 7530 8900
rect 7576 8888 7604 8919
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 8036 8965 8064 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11698 9024 11704 9036
rect 11348 8996 11704 9024
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7800 8928 8033 8956
rect 7800 8916 7806 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 8021 8919 8079 8925
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10778 8956 10784 8968
rect 10739 8928 10784 8956
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 11348 8965 11376 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 12250 8984 12256 9036
rect 12308 9024 12314 9036
rect 15473 9027 15531 9033
rect 12308 8996 14136 9024
rect 12308 8984 12314 8996
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11333 8919 11391 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12526 8956 12532 8968
rect 12207 8928 12532 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 14108 8965 14136 8996
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 16758 9024 16764 9036
rect 15519 8996 16764 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 18138 9024 18144 9036
rect 18051 8996 18144 9024
rect 18138 8984 18144 8996
rect 18196 9024 18202 9036
rect 19886 9024 19892 9036
rect 18196 8996 18368 9024
rect 18196 8984 18202 8996
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12768 8928 13001 8956
rect 12768 8916 12774 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 14424 8928 15761 8956
rect 14424 8916 14430 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 7524 8860 9045 8888
rect 7524 8848 7530 8860
rect 9033 8857 9045 8860
rect 9079 8857 9091 8891
rect 9033 8851 9091 8857
rect 10318 8848 10324 8900
rect 10376 8888 10382 8900
rect 10796 8888 10824 8916
rect 15764 8888 15792 8919
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15933 8959 15991 8965
rect 15933 8956 15945 8959
rect 15896 8928 15945 8956
rect 15896 8916 15902 8928
rect 15933 8925 15945 8928
rect 15979 8925 15991 8959
rect 16482 8956 16488 8968
rect 15933 8919 15991 8925
rect 16132 8928 16488 8956
rect 16022 8888 16028 8900
rect 10376 8860 12434 8888
rect 10376 8848 10382 8860
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 3602 8820 3608 8832
rect 2823 8792 3608 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 3881 8823 3939 8829
rect 3881 8820 3893 8823
rect 3844 8792 3893 8820
rect 3844 8780 3850 8792
rect 3881 8789 3893 8792
rect 3927 8789 3939 8823
rect 3881 8783 3939 8789
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4028 8792 4537 8820
rect 4028 8780 4034 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5721 8823 5779 8829
rect 5721 8820 5733 8823
rect 5408 8792 5733 8820
rect 5408 8780 5414 8792
rect 5721 8789 5733 8792
rect 5767 8789 5779 8823
rect 5721 8783 5779 8789
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8205 8823 8263 8829
rect 8205 8820 8217 8823
rect 8168 8792 8217 8820
rect 8168 8780 8174 8792
rect 8205 8789 8217 8792
rect 8251 8820 8263 8823
rect 10870 8820 10876 8832
rect 8251 8792 10876 8820
rect 8251 8789 8263 8792
rect 8205 8783 8263 8789
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 12406 8820 12434 8860
rect 14292 8860 15700 8888
rect 15764 8860 16028 8888
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 12406 8792 13185 8820
rect 13173 8789 13185 8792
rect 13219 8820 13231 8823
rect 13262 8820 13268 8832
rect 13219 8792 13268 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14090 8780 14096 8832
rect 14148 8820 14154 8832
rect 14292 8829 14320 8860
rect 14277 8823 14335 8829
rect 14277 8820 14289 8823
rect 14148 8792 14289 8820
rect 14148 8780 14154 8792
rect 14277 8789 14289 8792
rect 14323 8789 14335 8823
rect 14277 8783 14335 8789
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15286 8820 15292 8832
rect 15243 8792 15292 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15672 8820 15700 8860
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 16132 8820 16160 8928
rect 16482 8916 16488 8928
rect 16540 8956 16546 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16540 8928 16865 8956
rect 16540 8916 16546 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 17034 8956 17040 8968
rect 16995 8928 17040 8956
rect 16853 8919 16911 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 18049 8959 18107 8965
rect 17184 8928 17229 8956
rect 17184 8916 17190 8928
rect 18049 8925 18061 8959
rect 18095 8956 18107 8959
rect 18230 8956 18236 8968
rect 18095 8928 18236 8956
rect 18095 8925 18107 8928
rect 18049 8919 18107 8925
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 18340 8956 18368 8996
rect 19306 8996 19892 9024
rect 19306 8956 19334 8996
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 18340 8928 19334 8956
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 20533 8959 20591 8965
rect 20533 8956 20545 8959
rect 19760 8928 20545 8956
rect 19760 8916 19766 8928
rect 20533 8925 20545 8928
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 16669 8891 16727 8897
rect 16669 8857 16681 8891
rect 16715 8888 16727 8891
rect 19613 8891 19671 8897
rect 19613 8888 19625 8891
rect 16715 8860 19625 8888
rect 16715 8857 16727 8860
rect 16669 8851 16727 8857
rect 19613 8857 19625 8860
rect 19659 8857 19671 8891
rect 20714 8888 20720 8900
rect 20675 8860 20720 8888
rect 19613 8851 19671 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 15672 8792 16160 8820
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17589 8823 17647 8829
rect 17589 8820 17601 8823
rect 17552 8792 17601 8820
rect 17552 8780 17558 8792
rect 17589 8789 17601 8792
rect 17635 8789 17647 8823
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 17589 8783 17647 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 19518 8820 19524 8832
rect 19291 8792 19524 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 19794 8820 19800 8832
rect 19751 8792 19800 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 1104 8730 21436 8752
rect 1104 8678 7727 8730
rect 7779 8678 7791 8730
rect 7843 8678 7855 8730
rect 7907 8678 7919 8730
rect 7971 8678 7983 8730
rect 8035 8678 14504 8730
rect 14556 8678 14568 8730
rect 14620 8678 14632 8730
rect 14684 8678 14696 8730
rect 14748 8678 14760 8730
rect 14812 8678 21436 8730
rect 1104 8656 21436 8678
rect 2130 8616 2136 8628
rect 2091 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 2556 8588 3249 8616
rect 2556 8576 2562 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 4706 8616 4712 8628
rect 3237 8579 3295 8585
rect 3988 8588 4712 8616
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2148 8480 2176 8576
rect 2866 8548 2872 8560
rect 2779 8520 2872 8548
rect 2866 8508 2872 8520
rect 2924 8548 2930 8560
rect 3786 8548 3792 8560
rect 2924 8520 3792 8548
rect 2924 8508 2930 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 1903 8452 2176 8480
rect 2685 8483 2743 8489
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2774 8480 2780 8492
rect 2731 8452 2780 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3878 8480 3884 8492
rect 3099 8452 3884 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 1719 8384 2237 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2225 8381 2237 8384
rect 2271 8412 2283 8415
rect 2498 8412 2504 8424
rect 2271 8384 2504 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2976 8412 3004 8443
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 3988 8489 4016 8588
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8585 5043 8619
rect 5350 8616 5356 8628
rect 5311 8588 5356 8616
rect 4985 8579 5043 8585
rect 4246 8548 4252 8560
rect 4080 8520 4252 8548
rect 4080 8489 4108 8520
rect 4246 8508 4252 8520
rect 4304 8548 4310 8560
rect 5000 8548 5028 8579
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 6730 8616 6736 8628
rect 6691 8588 6736 8616
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 8812 8588 9321 8616
rect 8812 8576 8818 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 9416 8588 10916 8616
rect 4304 8520 5028 8548
rect 5445 8551 5503 8557
rect 4304 8508 4310 8520
rect 5445 8517 5457 8551
rect 5491 8548 5503 8551
rect 5534 8548 5540 8560
rect 5491 8520 5540 8548
rect 5491 8517 5503 8520
rect 5445 8511 5503 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 7650 8548 7656 8560
rect 7208 8520 7656 8548
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4341 8483 4399 8489
rect 4212 8452 4257 8480
rect 4212 8440 4218 8452
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 3142 8412 3148 8424
rect 2976 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3896 8412 3924 8440
rect 4350 8412 4378 8443
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 7208 8480 7236 8520
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 9416 8548 9444 8588
rect 8220 8520 9444 8548
rect 5040 8452 7236 8480
rect 7285 8483 7343 8489
rect 5040 8440 5046 8452
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7285 8443 7343 8449
rect 3896 8384 4378 8412
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5224 8384 5549 8412
rect 5224 8372 5230 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 7300 8412 7328 8443
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8110 8412 8116 8424
rect 6420 8384 7236 8412
rect 7300 8384 8116 8412
rect 6420 8372 6426 8384
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4062 8344 4068 8356
rect 3743 8316 4068 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 7208 8353 7236 8384
rect 7484 8356 7512 8384
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 4172 8316 7021 8344
rect 1946 8276 1952 8288
rect 1907 8248 1952 8276
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 3786 8236 3792 8288
rect 3844 8276 3850 8288
rect 4172 8276 4200 8316
rect 7009 8313 7021 8316
rect 7055 8313 7067 8347
rect 7009 8307 7067 8313
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8313 7251 8347
rect 7193 8307 7251 8313
rect 3844 8248 4200 8276
rect 3844 8236 3850 8248
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7116 8276 7144 8307
rect 7466 8304 7472 8356
rect 7524 8304 7530 8356
rect 8220 8276 8248 8520
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 9950 8548 9956 8560
rect 9548 8520 9628 8548
rect 9911 8520 9956 8548
rect 9548 8508 9554 8520
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8754 8480 8760 8492
rect 8527 8452 8760 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9600 8489 9628 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10888 8548 10916 8588
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 12069 8619 12127 8625
rect 11020 8588 11065 8616
rect 11020 8576 11026 8588
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 13906 8616 13912 8628
rect 12115 8588 13912 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 14056 8588 14197 8616
rect 14056 8576 14062 8588
rect 14185 8585 14197 8588
rect 14231 8616 14243 8619
rect 15102 8616 15108 8628
rect 14231 8588 15108 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 17954 8616 17960 8628
rect 16991 8588 17960 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 20257 8619 20315 8625
rect 20257 8616 20269 8619
rect 19208 8588 20269 8616
rect 19208 8576 19214 8588
rect 20257 8585 20269 8588
rect 20303 8585 20315 8619
rect 20257 8579 20315 8585
rect 14826 8548 14832 8560
rect 10888 8520 14832 8548
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 14918 8508 14924 8560
rect 14976 8548 14982 8560
rect 16390 8548 16396 8560
rect 14976 8520 16396 8548
rect 14976 8508 14982 8520
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 19429 8551 19487 8557
rect 19429 8548 19441 8551
rect 16908 8520 19441 8548
rect 16908 8508 16914 8520
rect 19429 8517 19441 8520
rect 19475 8517 19487 8551
rect 19429 8511 19487 8517
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9631 8452 9873 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8412 8355 8415
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8343 8384 8861 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9968 8412 9996 8508
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10778 8480 10784 8492
rect 10739 8452 10784 8480
rect 10505 8443 10563 8449
rect 9539 8384 9996 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 8864 8344 8892 8375
rect 10042 8344 10048 8356
rect 8864 8316 10048 8344
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10520 8344 10548 8443
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 13265 8483 13323 8489
rect 12492 8452 12537 8480
rect 12492 8440 12498 8452
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13722 8480 13728 8492
rect 13311 8452 13728 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 14182 8480 14188 8492
rect 14047 8452 14188 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 10686 8412 10692 8424
rect 10647 8384 10692 8412
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 11848 8384 12541 8412
rect 11848 8372 11854 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8412 12771 8415
rect 12802 8412 12808 8424
rect 12759 8384 12808 8412
rect 12759 8381 12771 8384
rect 12713 8375 12771 8381
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 14844 8412 14872 8508
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15470 8480 15476 8492
rect 15160 8452 15332 8480
rect 15431 8452 15476 8480
rect 15160 8440 15166 8452
rect 15194 8412 15200 8424
rect 14844 8384 15200 8412
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 14826 8344 14832 8356
rect 10520 8316 14832 8344
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 15102 8344 15108 8356
rect 15063 8316 15108 8344
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15304 8344 15332 8452
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 16114 8480 16120 8492
rect 15764 8452 16120 8480
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 15654 8412 15660 8424
rect 15611 8384 15660 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15764 8421 15792 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16482 8440 16488 8492
rect 16540 8480 16546 8492
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 16540 8452 17141 8480
rect 16540 8440 16546 8452
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18322 8480 18328 8492
rect 17911 8452 18328 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18690 8480 18696 8492
rect 18651 8452 18696 8480
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 19150 8480 19156 8492
rect 19111 8452 19156 8480
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 15896 8384 17417 8412
rect 15896 8372 15902 8384
rect 17405 8381 17417 8384
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 19352 8412 19380 8443
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 19576 8452 20177 8480
rect 19576 8440 19582 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 17644 8384 18552 8412
rect 17644 8372 17650 8384
rect 17034 8344 17040 8356
rect 15304 8316 17040 8344
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 18524 8353 18552 8384
rect 19168 8384 19380 8412
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 17184 8316 17969 8344
rect 17184 8304 17190 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 17957 8307 18015 8313
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8313 18567 8347
rect 18509 8307 18567 8313
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 19168 8344 19196 8384
rect 19705 8347 19763 8353
rect 19705 8344 19717 8347
rect 18656 8316 19196 8344
rect 19306 8316 19717 8344
rect 18656 8304 18662 8316
rect 6696 8248 8248 8276
rect 6696 8236 6702 8248
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 9364 8248 10517 8276
rect 9364 8236 9370 8248
rect 10505 8245 10517 8248
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 13354 8276 13360 8288
rect 11756 8248 13360 8276
rect 11756 8236 11762 8248
rect 13354 8236 13360 8248
rect 13412 8276 13418 8288
rect 13449 8279 13507 8285
rect 13449 8276 13461 8279
rect 13412 8248 13461 8276
rect 13412 8236 13418 8248
rect 13449 8245 13461 8248
rect 13495 8245 13507 8279
rect 13449 8239 13507 8245
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 16666 8276 16672 8288
rect 14976 8248 16672 8276
rect 14976 8236 14982 8248
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 17052 8276 17080 8304
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 17052 8248 17325 8276
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 19306 8276 19334 8316
rect 19705 8313 19717 8316
rect 19751 8313 19763 8347
rect 19705 8307 19763 8313
rect 19208 8248 19334 8276
rect 19208 8236 19214 8248
rect 1104 8186 21436 8208
rect 1104 8134 4338 8186
rect 4390 8134 4402 8186
rect 4454 8134 4466 8186
rect 4518 8134 4530 8186
rect 4582 8134 4594 8186
rect 4646 8134 11116 8186
rect 11168 8134 11180 8186
rect 11232 8134 11244 8186
rect 11296 8134 11308 8186
rect 11360 8134 11372 8186
rect 11424 8134 17893 8186
rect 17945 8134 17957 8186
rect 18009 8134 18021 8186
rect 18073 8134 18085 8186
rect 18137 8134 18149 8186
rect 18201 8134 21436 8186
rect 1104 8112 21436 8134
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9950 8072 9956 8084
rect 9180 8044 9956 8072
rect 9180 8032 9186 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 11900 8044 12388 8072
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 4982 8004 4988 8016
rect 1903 7976 4988 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 5442 8004 5448 8016
rect 5403 7976 5448 8004
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 9766 8004 9772 8016
rect 7760 7976 8064 8004
rect 9727 7976 9772 8004
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2188 7908 2636 7936
rect 2188 7896 2194 7908
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2608 7877 2636 7908
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 2832 7908 3832 7936
rect 2832 7896 2838 7908
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3804 7877 3832 7908
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4212 7908 4660 7936
rect 4212 7896 4218 7908
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7868 3847 7871
rect 3878 7868 3884 7880
rect 3835 7840 3884 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4632 7877 4660 7908
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5684 7908 5729 7936
rect 5828 7908 6224 7936
rect 5684 7896 5690 7908
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4028 7840 4445 7868
rect 4028 7828 4034 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 5316 7840 5365 7868
rect 5316 7828 5322 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5828 7868 5856 7908
rect 5353 7831 5411 7837
rect 5460 7840 5856 7868
rect 6089 7871 6147 7877
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 5460 7800 5488 7840
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 2004 7772 5488 7800
rect 2004 7760 2010 7772
rect 2314 7732 2320 7744
rect 2275 7704 2320 7732
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 3752 7704 4537 7732
rect 3752 7692 3758 7704
rect 4525 7701 4537 7704
rect 4571 7701 4583 7735
rect 4525 7695 4583 7701
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 6104 7732 6132 7831
rect 6196 7800 6224 7908
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 7760 7936 7788 7976
rect 6788 7908 7788 7936
rect 6788 7896 6794 7908
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8036 7936 8064 7976
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10134 7964 10140 8016
rect 10192 8004 10198 8016
rect 11900 8013 11928 8044
rect 11885 8007 11943 8013
rect 10192 7976 11836 8004
rect 10192 7964 10198 7976
rect 10226 7936 10232 7948
rect 7892 7908 7972 7936
rect 8036 7908 10232 7936
rect 7892 7896 7898 7908
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7432 7840 7665 7868
rect 7432 7828 7438 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7944 7868 7972 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11698 7936 11704 7948
rect 10428 7908 11704 7936
rect 8570 7868 8576 7880
rect 7944 7840 8576 7868
rect 7653 7831 7711 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 9088 7840 9137 7868
rect 9088 7828 9094 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9582 7868 9588 7880
rect 9543 7840 9588 7868
rect 9125 7831 9183 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9732 7840 9781 7868
rect 9732 7828 9738 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10318 7868 10324 7880
rect 10091 7840 10324 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10428 7877 10456 7908
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 10870 7868 10876 7880
rect 10643 7840 10876 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11238 7868 11244 7880
rect 11199 7840 11244 7868
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11808 7868 11836 7976
rect 11885 7973 11897 8007
rect 11931 7973 11943 8007
rect 12360 8004 12388 8044
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12492 8044 12909 8072
rect 12492 8032 12498 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 13354 8072 13360 8084
rect 13315 8044 13360 8072
rect 12897 8035 12955 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 15470 8072 15476 8084
rect 15335 8044 15476 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16666 8072 16672 8084
rect 15712 8044 16672 8072
rect 15712 8032 15718 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16816 8044 16957 8072
rect 16816 8032 16822 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 19426 8072 19432 8084
rect 16945 8035 17003 8041
rect 17052 8044 19432 8072
rect 12802 8004 12808 8016
rect 12360 7976 12808 8004
rect 11885 7967 11943 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 14737 8007 14795 8013
rect 14737 7973 14749 8007
rect 14783 8004 14795 8007
rect 15930 8004 15936 8016
rect 14783 7976 15936 8004
rect 14783 7973 14795 7976
rect 14737 7967 14795 7973
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 16114 7964 16120 8016
rect 16172 8004 16178 8016
rect 17052 8004 17080 8044
rect 19426 8032 19432 8044
rect 19484 8072 19490 8084
rect 20254 8072 20260 8084
rect 19484 8044 20260 8072
rect 19484 8032 19490 8044
rect 20254 8032 20260 8044
rect 20312 8032 20318 8084
rect 16172 7976 17080 8004
rect 16172 7964 16178 7976
rect 17494 7964 17500 8016
rect 17552 8004 17558 8016
rect 18322 8004 18328 8016
rect 17552 7976 18328 8004
rect 17552 7964 17558 7976
rect 18322 7964 18328 7976
rect 18380 7964 18386 8016
rect 19518 8004 19524 8016
rect 18432 7976 19524 8004
rect 11974 7936 11980 7948
rect 11887 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7936 12038 7948
rect 15749 7939 15807 7945
rect 12032 7908 13124 7936
rect 12032 7896 12038 7908
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11808 7840 12081 7868
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7868 12219 7871
rect 12250 7868 12256 7880
rect 12207 7840 12256 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12618 7868 12624 7880
rect 12483 7840 12624 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 6196 7772 7757 7800
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 7745 7763 7803 7769
rect 8846 7760 8852 7812
rect 8904 7800 8910 7812
rect 8904 7772 11652 7800
rect 8904 7760 8910 7772
rect 5500 7704 6132 7732
rect 5500 7692 5506 7704
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 6236 7704 6285 7732
rect 6236 7692 6242 7704
rect 6273 7701 6285 7704
rect 6319 7701 6331 7735
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 6273 7695 6331 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 10502 7732 10508 7744
rect 8987 7704 10508 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11146 7732 11152 7744
rect 11103 7704 11152 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11624 7732 11652 7772
rect 11698 7760 11704 7812
rect 11756 7800 11762 7812
rect 12360 7800 12388 7831
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13096 7877 13124 7908
rect 15396 7908 15608 7936
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12860 7840 12909 7868
rect 12860 7828 12866 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7868 13231 7871
rect 13262 7868 13268 7880
rect 13219 7840 13268 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 11756 7772 12388 7800
rect 11756 7760 11762 7772
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13464 7800 13492 7831
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 13964 7840 14565 7868
rect 13964 7828 13970 7840
rect 14553 7837 14565 7840
rect 14599 7868 14611 7871
rect 15010 7868 15016 7880
rect 14599 7840 15016 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 12584 7772 13492 7800
rect 12584 7760 12590 7772
rect 13722 7732 13728 7744
rect 11624 7704 13728 7732
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15396 7732 15424 7908
rect 15580 7877 15608 7908
rect 15749 7905 15761 7939
rect 15795 7936 15807 7939
rect 16298 7936 16304 7948
rect 15795 7908 16304 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 17862 7936 17868 7948
rect 16816 7908 17868 7936
rect 16816 7896 16822 7908
rect 17862 7896 17868 7908
rect 17920 7936 17926 7948
rect 18432 7936 18460 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 17920 7908 18460 7936
rect 17920 7896 17926 7908
rect 15473 7871 15531 7877
rect 15473 7837 15485 7871
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7837 15623 7871
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15565 7831 15623 7837
rect 15488 7800 15516 7831
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 15948 7840 16865 7868
rect 15948 7800 15976 7840
rect 16853 7837 16865 7840
rect 16899 7868 16911 7871
rect 17034 7868 17040 7880
rect 16899 7840 17040 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17494 7868 17500 7880
rect 17455 7840 17500 7868
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 18230 7868 18236 7880
rect 17635 7840 18236 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 18230 7828 18236 7840
rect 18288 7868 18294 7880
rect 18432 7877 18460 7908
rect 19444 7908 19901 7936
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 18288 7840 18337 7868
rect 18288 7828 18294 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18598 7868 18604 7880
rect 18559 7840 18604 7868
rect 18417 7831 18475 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7868 18751 7871
rect 18782 7868 18788 7880
rect 18739 7840 18788 7868
rect 18739 7837 18751 7840
rect 18693 7831 18751 7837
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19444 7877 19472 7908
rect 19889 7905 19901 7908
rect 19935 7905 19947 7939
rect 19889 7899 19947 7905
rect 19426 7871 19484 7877
rect 19426 7868 19438 7871
rect 19116 7840 19438 7868
rect 19116 7828 19122 7840
rect 19426 7837 19438 7840
rect 19472 7837 19484 7871
rect 19426 7831 19484 7837
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 15488 7772 15976 7800
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 19812 7800 19840 7831
rect 20530 7800 20536 7812
rect 16724 7772 19288 7800
rect 16724 7760 16730 7772
rect 15470 7732 15476 7744
rect 15396 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 17954 7732 17960 7744
rect 15804 7704 17960 7732
rect 15804 7692 15810 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18506 7732 18512 7744
rect 18187 7704 18512 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 18966 7732 18972 7744
rect 18656 7704 18972 7732
rect 18656 7692 18662 7704
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 19260 7741 19288 7772
rect 19444 7772 19840 7800
rect 20491 7772 20536 7800
rect 19245 7735 19303 7741
rect 19245 7701 19257 7735
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19444 7741 19472 7772
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19392 7704 19441 7732
rect 19392 7692 19398 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 20622 7732 20628 7744
rect 20583 7704 20628 7732
rect 19429 7695 19487 7701
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 1104 7642 21436 7664
rect 1104 7590 7727 7642
rect 7779 7590 7791 7642
rect 7843 7590 7855 7642
rect 7907 7590 7919 7642
rect 7971 7590 7983 7642
rect 8035 7590 14504 7642
rect 14556 7590 14568 7642
rect 14620 7590 14632 7642
rect 14684 7590 14696 7642
rect 14748 7590 14760 7642
rect 14812 7590 21436 7642
rect 1104 7568 21436 7590
rect 6730 7528 6736 7540
rect 2746 7500 6736 7528
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 2746 7256 2774 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7466 7528 7472 7540
rect 7055 7500 7472 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7497 8539 7531
rect 8481 7491 8539 7497
rect 2976 7432 4200 7460
rect 2976 7401 3004 7432
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 3694 7392 3700 7404
rect 3655 7364 3700 7392
rect 2961 7355 3019 7361
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 4172 7401 4200 7432
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 6546 7460 6552 7472
rect 5316 7432 6552 7460
rect 5316 7420 5322 7432
rect 6546 7420 6552 7432
rect 6604 7460 6610 7472
rect 8496 7460 8524 7491
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 9640 7500 9689 7528
rect 9640 7488 9646 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 10134 7528 10140 7540
rect 9907 7500 10140 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 10744 7500 11989 7528
rect 10744 7488 10750 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 11977 7491 12035 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 13630 7528 13636 7540
rect 12308 7500 12388 7528
rect 13591 7500 13636 7528
rect 12308 7488 12314 7500
rect 10778 7460 10784 7472
rect 6604 7432 7144 7460
rect 8496 7432 10784 7460
rect 6604 7420 6610 7432
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3844 7364 3893 7392
rect 3844 7352 3850 7364
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4246 7392 4252 7404
rect 4203 7364 4252 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4706 7392 4712 7404
rect 4387 7364 4712 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4706 7352 4712 7364
rect 4764 7392 4770 7404
rect 5350 7392 5356 7404
rect 4764 7364 5356 7392
rect 4764 7352 4770 7364
rect 5350 7352 5356 7364
rect 5408 7392 5414 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5408 7364 5457 7392
rect 5408 7352 5414 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 6362 7392 6368 7404
rect 5960 7364 6368 7392
rect 5960 7352 5966 7364
rect 6362 7352 6368 7364
rect 6420 7392 6426 7404
rect 7116 7401 7144 7432
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 6825 7396 6883 7401
rect 6656 7395 6883 7396
rect 6656 7392 6837 7395
rect 6420 7368 6837 7392
rect 6420 7364 6684 7368
rect 6420 7352 6426 7364
rect 6825 7361 6837 7368
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8294 7392 8300 7404
rect 8255 7364 8300 7392
rect 8021 7355 8079 7361
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 2087 7228 2774 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 3988 7256 4016 7287
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 8036 7324 8064 7355
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8812 7364 8953 7392
rect 8812 7352 8818 7364
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 9950 7392 9956 7404
rect 9640 7364 9956 7392
rect 9640 7352 9646 7364
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10594 7392 10600 7404
rect 10275 7364 10600 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11238 7392 11244 7404
rect 11011 7364 11244 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11793 7395 11851 7401
rect 11563 7364 11744 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 4948 7296 8064 7324
rect 4948 7284 4954 7296
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8168 7296 8213 7324
rect 8168 7284 8174 7296
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9732 7296 9781 7324
rect 9732 7284 9738 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 3936 7228 4016 7256
rect 3936 7216 3942 7228
rect 4154 7216 4160 7268
rect 4212 7256 4218 7268
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 4212 7228 5549 7256
rect 4212 7216 4218 7228
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 6641 7259 6699 7265
rect 6641 7256 6653 7259
rect 5583 7228 6653 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 6641 7225 6653 7228
rect 6687 7225 6699 7259
rect 9784 7256 9812 7287
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 10468 7296 11621 7324
rect 10468 7284 10474 7296
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 10226 7256 10232 7268
rect 9784 7228 10232 7256
rect 6641 7219 6699 7225
rect 10226 7216 10232 7228
rect 10284 7256 10290 7268
rect 11716 7256 11744 7364
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11974 7392 11980 7404
rect 11839 7364 11980 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7392 12038 7404
rect 12250 7392 12256 7404
rect 12032 7364 12256 7392
rect 12032 7352 12038 7364
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12360 7324 12388 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 17920 7500 18276 7528
rect 17920 7488 17926 7500
rect 18248 7469 18276 7500
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 18601 7531 18659 7537
rect 18601 7497 18613 7531
rect 18647 7528 18659 7531
rect 18647 7500 19104 7528
rect 18647 7497 18659 7500
rect 18601 7491 18659 7497
rect 13449 7463 13507 7469
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 15381 7463 15439 7469
rect 13495 7432 13676 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 12710 7392 12716 7404
rect 12671 7364 12716 7392
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13538 7392 13544 7404
rect 13499 7364 13544 7392
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13648 7392 13676 7432
rect 15381 7429 15393 7463
rect 15427 7460 15439 7463
rect 18233 7463 18291 7469
rect 15427 7432 16712 7460
rect 15427 7429 15439 7432
rect 15381 7423 15439 7429
rect 13814 7392 13820 7404
rect 13648 7364 13820 7392
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13964 7364 14013 7392
rect 13964 7352 13970 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14918 7392 14924 7404
rect 14879 7364 14924 7392
rect 14001 7355 14059 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 16022 7401 16028 7404
rect 15979 7395 16028 7401
rect 15528 7364 15884 7392
rect 15528 7352 15534 7364
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 12360 7296 13737 7324
rect 13725 7293 13737 7296
rect 13771 7324 13783 7327
rect 15102 7324 15108 7336
rect 13771 7296 15108 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 15252 7296 15761 7324
rect 15252 7284 15258 7296
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15856 7324 15884 7364
rect 15979 7361 15991 7395
rect 16025 7361 16028 7395
rect 15979 7355 16028 7361
rect 16022 7352 16028 7355
rect 16080 7352 16086 7404
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16482 7392 16488 7404
rect 16163 7364 16488 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16684 7401 16712 7432
rect 18233 7429 18245 7463
rect 18279 7429 18291 7463
rect 18340 7460 18368 7488
rect 19076 7472 19104 7500
rect 19058 7460 19064 7472
rect 18340 7432 18460 7460
rect 19019 7432 19064 7460
rect 18233 7423 18291 7429
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 16669 7355 16727 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17003 7395 17061 7401
rect 17003 7361 17015 7395
rect 17049 7392 17061 7395
rect 17049 7361 17080 7392
rect 17003 7355 17080 7361
rect 17052 7324 17080 7355
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 17184 7364 17233 7392
rect 17184 7352 17190 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7392 18107 7395
rect 18138 7392 18144 7404
rect 18095 7364 18144 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18322 7392 18328 7404
rect 18283 7364 18328 7392
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18432 7401 18460 7432
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 18874 7392 18880 7404
rect 18656 7364 18880 7392
rect 18656 7352 18662 7364
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 19208 7364 19257 7392
rect 19208 7352 19214 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 20349 7395 20407 7401
rect 20349 7392 20361 7395
rect 19245 7355 19303 7361
rect 19352 7364 20361 7392
rect 19352 7324 19380 7364
rect 20349 7361 20361 7364
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 15856 7296 16068 7324
rect 15749 7287 15807 7293
rect 13538 7256 13544 7268
rect 10284 7228 11744 7256
rect 11808 7228 13544 7256
rect 10284 7216 10290 7228
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3970 7188 3976 7200
rect 3099 7160 3976 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 6052 7160 6377 7188
rect 6052 7148 6058 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6730 7188 6736 7200
rect 6691 7160 6736 7188
rect 6365 7151 6423 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7248 7160 8033 7188
rect 7248 7148 7254 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 9125 7191 9183 7197
rect 9125 7157 9137 7191
rect 9171 7188 9183 7191
rect 9306 7188 9312 7200
rect 9171 7160 9312 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 10134 7188 10140 7200
rect 10095 7160 10140 7188
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11808 7197 11836 7228
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 15436 7228 15853 7256
rect 15436 7216 15442 7228
rect 15764 7200 15792 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 16040 7256 16068 7296
rect 16960 7296 17080 7324
rect 18524 7296 19380 7324
rect 16960 7256 16988 7296
rect 16040 7228 16988 7256
rect 17037 7259 17095 7265
rect 15841 7219 15899 7225
rect 17037 7225 17049 7259
rect 17083 7256 17095 7259
rect 17083 7228 18184 7256
rect 17083 7225 17095 7228
rect 17037 7219 17095 7225
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7157 11851 7191
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 11793 7151 11851 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13780 7160 13921 7188
rect 13780 7148 13786 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 13909 7151 13967 7157
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15286 7188 15292 7200
rect 14783 7160 15292 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7148 15810 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 16356 7160 17141 7188
rect 16356 7148 16362 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 18156 7188 18184 7228
rect 18524 7188 18552 7296
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 20220 7296 20453 7324
rect 20220 7284 20226 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 20548 7256 20576 7287
rect 20312 7228 20576 7256
rect 20312 7216 20318 7228
rect 18156 7160 18552 7188
rect 17129 7151 17187 7157
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 18656 7160 19441 7188
rect 18656 7148 18662 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19944 7160 19993 7188
rect 19944 7148 19950 7160
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 1104 7098 21436 7120
rect 1104 7046 4338 7098
rect 4390 7046 4402 7098
rect 4454 7046 4466 7098
rect 4518 7046 4530 7098
rect 4582 7046 4594 7098
rect 4646 7046 11116 7098
rect 11168 7046 11180 7098
rect 11232 7046 11244 7098
rect 11296 7046 11308 7098
rect 11360 7046 11372 7098
rect 11424 7046 17893 7098
rect 17945 7046 17957 7098
rect 18009 7046 18021 7098
rect 18073 7046 18085 7098
rect 18137 7046 18149 7098
rect 18201 7046 21436 7098
rect 1104 7024 21436 7046
rect 2866 6984 2872 6996
rect 2779 6956 2872 6984
rect 2866 6944 2872 6956
rect 2924 6984 2930 6996
rect 3786 6984 3792 6996
rect 2924 6956 3792 6984
rect 2924 6944 2930 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4304 6956 4752 6984
rect 4304 6944 4310 6956
rect 4724 6916 4752 6956
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 8294 6984 8300 6996
rect 5408 6956 8300 6984
rect 5408 6944 5414 6956
rect 5997 6919 6055 6925
rect 5997 6916 6009 6919
rect 4724 6888 6009 6916
rect 5997 6885 6009 6888
rect 6043 6885 6055 6919
rect 5997 6879 6055 6885
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 3510 6848 3516 6860
rect 2271 6820 3516 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 4246 6848 4252 6860
rect 3712 6820 4252 6848
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2372 6752 2789 6780
rect 2372 6740 2378 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 1949 6715 2007 6721
rect 1949 6681 1961 6715
rect 1995 6712 2007 6715
rect 3712 6712 3740 6820
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 3844 6752 3889 6780
rect 3844 6740 3850 6752
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 4028 6752 4077 6780
rect 4028 6740 4034 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 5350 6780 5356 6792
rect 5311 6752 5356 6780
rect 4525 6743 4583 6749
rect 4540 6712 4568 6743
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6196 6789 6224 6956
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 10686 6984 10692 6996
rect 10192 6956 10692 6984
rect 10192 6944 10198 6956
rect 10686 6944 10692 6956
rect 10744 6984 10750 6996
rect 12158 6984 12164 6996
rect 10744 6956 12164 6984
rect 10744 6944 10750 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 16022 6984 16028 6996
rect 15212 6956 16028 6984
rect 6914 6916 6920 6928
rect 6380 6888 6920 6916
rect 6380 6848 6408 6888
rect 6914 6876 6920 6888
rect 6972 6876 6978 6928
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7837 6919 7895 6925
rect 7837 6916 7849 6919
rect 7340 6888 7849 6916
rect 7340 6876 7346 6888
rect 7837 6885 7849 6888
rect 7883 6885 7895 6919
rect 8110 6916 8116 6928
rect 7837 6879 7895 6885
rect 7944 6888 8116 6916
rect 6288 6820 6408 6848
rect 6457 6851 6515 6857
rect 6288 6789 6316 6820
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 7098 6848 7104 6860
rect 6503 6820 7104 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 7944 6857 7972 6888
rect 8110 6876 8116 6888
rect 8168 6916 8174 6928
rect 14366 6916 14372 6928
rect 8168 6888 14372 6916
rect 8168 6876 8174 6888
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 15212 6916 15240 6956
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 18414 6984 18420 6996
rect 16540 6956 18420 6984
rect 16540 6944 16546 6956
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 18601 6987 18659 6993
rect 18601 6953 18613 6987
rect 18647 6984 18659 6987
rect 18782 6984 18788 6996
rect 18647 6956 18788 6984
rect 18647 6953 18659 6956
rect 18601 6947 18659 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 20162 6984 20168 6996
rect 20123 6956 20168 6984
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 14936 6888 15240 6916
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7708 6820 7941 6848
rect 7708 6808 7714 6820
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7929 6811 7987 6817
rect 8036 6820 8217 6848
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6273 6743 6331 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 1995 6684 3740 6712
rect 3896 6684 4568 6712
rect 5368 6712 5396 6740
rect 7208 6712 7236 6743
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 8036 6780 8064 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8386 6848 8392 6860
rect 8347 6820 8392 6848
rect 8205 6811 8263 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9582 6848 9588 6860
rect 8772 6820 9588 6848
rect 7432 6752 8064 6780
rect 8113 6783 8171 6789
rect 7432 6740 7438 6752
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8772 6780 8800 6820
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10468 6820 11069 6848
rect 10468 6808 10474 6820
rect 11057 6817 11069 6820
rect 11103 6848 11115 6851
rect 11606 6848 11612 6860
rect 11103 6820 11612 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 14936 6857 14964 6888
rect 15654 6876 15660 6928
rect 15712 6916 15718 6928
rect 17589 6919 17647 6925
rect 17589 6916 17601 6919
rect 15712 6888 17601 6916
rect 15712 6876 15718 6888
rect 17589 6885 17601 6888
rect 17635 6916 17647 6919
rect 18690 6916 18696 6928
rect 17635 6888 18696 6916
rect 17635 6885 17647 6888
rect 17589 6879 17647 6885
rect 18690 6876 18696 6888
rect 18748 6876 18754 6928
rect 19150 6876 19156 6928
rect 19208 6916 19214 6928
rect 19208 6888 19472 6916
rect 19208 6876 19214 6888
rect 12805 6851 12863 6857
rect 12805 6848 12817 6851
rect 12032 6820 12817 6848
rect 12032 6808 12038 6820
rect 12805 6817 12817 6820
rect 12851 6817 12863 6851
rect 12805 6811 12863 6817
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6817 14979 6851
rect 14921 6811 14979 6817
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15068 6820 15393 6848
rect 15068 6808 15074 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 17034 6848 17040 6860
rect 16071 6820 17040 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 19334 6848 19340 6860
rect 18187 6820 19340 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 19444 6848 19472 6888
rect 19889 6851 19947 6857
rect 19889 6848 19901 6851
rect 19444 6820 19901 6848
rect 19889 6817 19901 6820
rect 19935 6848 19947 6851
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 19935 6820 20453 6848
rect 19935 6817 19947 6820
rect 19889 6811 19947 6817
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 8938 6780 8944 6792
rect 8159 6752 8800 6780
rect 8899 6752 8944 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9272 6752 9781 6780
rect 9272 6740 9278 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6749 10839 6783
rect 10962 6780 10968 6792
rect 10923 6752 10968 6780
rect 10781 6743 10839 6749
rect 8386 6712 8392 6724
rect 5368 6684 8392 6712
rect 1995 6681 2007 6684
rect 1949 6675 2007 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2096 6616 2141 6644
rect 2096 6604 2102 6616
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3896 6653 3924 6684
rect 8386 6672 8392 6684
rect 8444 6672 8450 6724
rect 9582 6712 9588 6724
rect 8956 6684 9444 6712
rect 9543 6684 9588 6712
rect 3887 6647 3945 6653
rect 3887 6644 3899 6647
rect 2648 6616 3899 6644
rect 2648 6604 2654 6616
rect 3887 6613 3899 6616
rect 3933 6613 3945 6647
rect 3887 6607 3945 6613
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4154 6644 4160 6656
rect 4019 6616 4160 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4614 6644 4620 6656
rect 4575 6616 4620 6644
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 7009 6647 7067 6653
rect 7009 6644 7021 6647
rect 5592 6616 7021 6644
rect 5592 6604 5598 6616
rect 7009 6613 7021 6616
rect 7055 6613 7067 6647
rect 7009 6607 7067 6613
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 8956 6644 8984 6684
rect 9122 6644 9128 6656
rect 8067 6616 8984 6644
rect 9083 6616 9128 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9416 6644 9444 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9858 6712 9864 6724
rect 9771 6684 9864 6712
rect 9784 6644 9812 6684
rect 9858 6672 9864 6684
rect 9916 6712 9922 6724
rect 10796 6712 10824 6743
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11756 6752 11897 6780
rect 11756 6740 11762 6752
rect 11885 6749 11897 6752
rect 11931 6780 11943 6783
rect 12526 6780 12532 6792
rect 11931 6752 12434 6780
rect 12487 6752 12532 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12406 6724 12434 6752
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 12621 6743 12679 6749
rect 11606 6712 11612 6724
rect 9916 6684 10732 6712
rect 10796 6684 11612 6712
rect 9916 6672 9922 6684
rect 9950 6644 9956 6656
rect 9416 6616 9812 6644
rect 9911 6616 9956 6644
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10704 6644 10732 6684
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 12158 6712 12164 6724
rect 11716 6684 12164 6712
rect 11716 6644 11744 6684
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 12406 6684 12440 6724
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 10704 6616 11744 6644
rect 11977 6647 12035 6653
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12544 6644 12572 6740
rect 12636 6712 12664 6743
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 13780 6752 14197 6780
rect 13780 6740 13786 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 15102 6780 15108 6792
rect 15063 6752 15108 6780
rect 14185 6743 14243 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 15654 6780 15660 6792
rect 15335 6752 15660 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 16117 6783 16175 6789
rect 16117 6782 16129 6783
rect 15994 6780 16129 6782
rect 15804 6754 16129 6780
rect 15804 6752 16022 6754
rect 15804 6740 15810 6752
rect 16117 6749 16129 6754
rect 16163 6749 16175 6783
rect 16758 6780 16764 6792
rect 16719 6752 16764 6780
rect 16117 6743 16175 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 16908 6752 17509 6780
rect 16908 6740 16914 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 12636 6684 13369 6712
rect 13357 6681 13369 6684
rect 13403 6712 13415 6715
rect 13446 6712 13452 6724
rect 13403 6684 13452 6712
rect 13403 6681 13415 6684
rect 13357 6675 13415 6681
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 15841 6715 15899 6721
rect 14884 6684 15240 6712
rect 14884 6672 14890 6684
rect 12023 6616 12572 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12768 6616 12817 6644
rect 12768 6604 12774 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14366 6644 14372 6656
rect 14323 6616 14372 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14918 6644 14924 6656
rect 14879 6616 14924 6644
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 15212 6644 15240 6684
rect 15841 6681 15853 6715
rect 15887 6712 15899 6715
rect 16868 6712 16896 6740
rect 15887 6684 16896 6712
rect 18340 6712 18368 6743
rect 18414 6740 18420 6792
rect 18472 6780 18478 6792
rect 18690 6780 18696 6792
rect 18472 6752 18517 6780
rect 18651 6752 18696 6780
rect 18472 6740 18478 6752
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19116 6752 19257 6780
rect 19116 6740 19122 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 20070 6780 20076 6792
rect 19475 6752 19564 6780
rect 20031 6752 20076 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19150 6712 19156 6724
rect 18340 6684 19156 6712
rect 15887 6681 15899 6684
rect 15841 6675 15899 6681
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 19536 6712 19564 6752
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 19260 6684 19564 6712
rect 20088 6712 20116 6740
rect 20349 6715 20407 6721
rect 20349 6712 20361 6715
rect 20088 6684 20361 6712
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 15068 6616 15113 6644
rect 15212 6616 16313 6644
rect 15068 6604 15074 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16850 6644 16856 6656
rect 16811 6616 16856 6644
rect 16301 6607 16359 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18322 6644 18328 6656
rect 18012 6616 18328 6644
rect 18012 6604 18018 6616
rect 18322 6604 18328 6616
rect 18380 6644 18386 6656
rect 19260 6644 19288 6684
rect 19426 6644 19432 6656
rect 18380 6616 19288 6644
rect 19387 6616 19432 6644
rect 18380 6604 18386 6616
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 19536 6644 19564 6684
rect 20349 6681 20361 6684
rect 20395 6681 20407 6715
rect 20349 6675 20407 6681
rect 20622 6644 20628 6656
rect 19536 6616 20628 6644
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 1104 6554 21436 6576
rect 1104 6502 7727 6554
rect 7779 6502 7791 6554
rect 7843 6502 7855 6554
rect 7907 6502 7919 6554
rect 7971 6502 7983 6554
rect 8035 6502 14504 6554
rect 14556 6502 14568 6554
rect 14620 6502 14632 6554
rect 14684 6502 14696 6554
rect 14748 6502 14760 6554
rect 14812 6502 21436 6554
rect 1104 6480 21436 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 5166 6440 5172 6452
rect 3200 6412 5172 6440
rect 3200 6400 3206 6412
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 7374 6440 7380 6452
rect 6512 6412 7380 6440
rect 6512 6400 6518 6412
rect 7374 6400 7380 6412
rect 7432 6440 7438 6452
rect 9490 6440 9496 6452
rect 7432 6412 7512 6440
rect 9451 6412 9496 6440
rect 7432 6400 7438 6412
rect 2498 6332 2504 6384
rect 2556 6372 2562 6384
rect 3329 6375 3387 6381
rect 3329 6372 3341 6375
rect 2556 6344 3341 6372
rect 2556 6332 2562 6344
rect 3329 6341 3341 6344
rect 3375 6341 3387 6375
rect 4614 6372 4620 6384
rect 3329 6335 3387 6341
rect 3436 6344 4620 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1762 6304 1768 6316
rect 1627 6276 1768 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2240 6236 2268 6267
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2590 6304 2596 6316
rect 2372 6276 2417 6304
rect 2551 6276 2596 6304
rect 2372 6264 2378 6276
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 3016 6276 3065 6304
rect 3016 6264 3022 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3436 6304 3464 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 3191 6276 3464 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 2501 6239 2559 6245
rect 2240 6208 2360 6236
rect 2332 6168 2360 6208
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2866 6236 2872 6248
rect 2547 6208 2872 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3160 6236 3188 6267
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3844 6276 3985 6304
rect 3844 6264 3850 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4433 6307 4491 6313
rect 4120 6276 4165 6304
rect 4120 6264 4126 6276
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4706 6304 4712 6316
rect 4479 6276 4712 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4706 6264 4712 6276
rect 4764 6304 4770 6316
rect 4890 6304 4896 6316
rect 4764 6276 4896 6304
rect 4764 6264 4770 6276
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 5040 6276 5089 6304
rect 5040 6264 5046 6276
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7190 6304 7196 6316
rect 6687 6276 7196 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7190 6264 7196 6276
rect 7248 6304 7254 6316
rect 7385 6307 7443 6313
rect 7248 6276 7328 6304
rect 7248 6264 7254 6276
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 2976 6208 3188 6236
rect 3252 6208 4169 6236
rect 2976 6180 3004 6208
rect 2958 6168 2964 6180
rect 2332 6140 2964 6168
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3053 6171 3111 6177
rect 3053 6137 3065 6171
rect 3099 6168 3111 6171
rect 3252 6168 3280 6208
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4798 6236 4804 6248
rect 4295 6208 4804 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7300 6236 7328 6276
rect 7385 6273 7397 6307
rect 7431 6304 7443 6307
rect 7484 6304 7512 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9950 6440 9956 6452
rect 9911 6412 9956 6440
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10870 6440 10876 6452
rect 10831 6412 10876 6440
rect 10870 6400 10876 6412
rect 10928 6440 10934 6452
rect 10928 6412 12020 6440
rect 10928 6400 10934 6412
rect 9858 6372 9864 6384
rect 9771 6344 9864 6372
rect 9858 6332 9864 6344
rect 9916 6372 9922 6384
rect 10594 6372 10600 6384
rect 9916 6344 10600 6372
rect 9916 6332 9922 6344
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 10888 6344 11928 6372
rect 8386 6304 8392 6316
rect 7431 6276 7512 6304
rect 8347 6276 8392 6304
rect 7431 6273 7443 6276
rect 7385 6267 7443 6273
rect 8386 6264 8392 6276
rect 8444 6304 8450 6316
rect 9030 6304 9036 6316
rect 8444 6276 9036 6304
rect 8444 6264 8450 6276
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9140 6276 10640 6304
rect 9140 6236 9168 6276
rect 6972 6208 7017 6236
rect 7300 6208 9168 6236
rect 10137 6239 10195 6245
rect 6972 6196 6978 6208
rect 10137 6205 10149 6239
rect 10183 6205 10195 6239
rect 10612 6236 10640 6276
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10744 6276 10793 6304
rect 10744 6264 10750 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 10888 6236 10916 6344
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11664 6276 11713 6304
rect 11664 6264 11670 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 10612 6208 10916 6236
rect 10137 6199 10195 6205
rect 3099 6140 3280 6168
rect 3099 6137 3111 6140
rect 3053 6131 3111 6137
rect 6086 6128 6092 6180
rect 6144 6168 6150 6180
rect 8205 6171 8263 6177
rect 6144 6140 6776 6168
rect 6144 6128 6150 6140
rect 6748 6112 6776 6140
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 10152 6168 10180 6199
rect 10962 6196 10968 6248
rect 11020 6236 11026 6248
rect 11900 6236 11928 6344
rect 11992 6313 12020 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 15010 6440 15016 6452
rect 12216 6412 15016 6440
rect 12216 6400 12222 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 19794 6440 19800 6452
rect 15120 6412 17816 6440
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12621 6375 12679 6381
rect 12621 6372 12633 6375
rect 12400 6344 12633 6372
rect 12400 6332 12406 6344
rect 12621 6341 12633 6344
rect 12667 6341 12679 6375
rect 12621 6335 12679 6341
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 14553 6375 14611 6381
rect 14553 6372 14565 6375
rect 13320 6344 14565 6372
rect 13320 6332 13326 6344
rect 14553 6341 14565 6344
rect 14599 6341 14611 6375
rect 14553 6335 14611 6341
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 15120 6372 15148 6412
rect 16022 6372 16028 6384
rect 14700 6344 15148 6372
rect 15764 6344 16028 6372
rect 14700 6332 14706 6344
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 13280 6304 13308 6332
rect 13446 6304 13452 6316
rect 12483 6276 13308 6304
rect 13407 6276 13452 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13630 6304 13636 6316
rect 13591 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13771 6276 14197 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14185 6273 14197 6276
rect 14231 6304 14243 6307
rect 14274 6304 14280 6316
rect 14231 6276 14280 6304
rect 14231 6273 14243 6276
rect 14185 6267 14243 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 13262 6236 13268 6248
rect 11020 6208 11652 6236
rect 11900 6208 13268 6236
rect 11020 6196 11026 6208
rect 10594 6168 10600 6180
rect 8251 6140 9674 6168
rect 10152 6140 10600 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 2130 6100 2136 6112
rect 1443 6072 2136 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4212 6072 4905 6100
rect 4212 6060 4218 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 6328 6072 6469 6100
rect 6328 6060 6334 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6788 6072 6837 6100
rect 6788 6060 6794 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7374 6100 7380 6112
rect 6972 6072 7380 6100
rect 6972 6060 6978 6072
rect 7374 6060 7380 6072
rect 7432 6100 7438 6112
rect 7469 6103 7527 6109
rect 7469 6100 7481 6103
rect 7432 6072 7481 6100
rect 7432 6060 7438 6072
rect 7469 6069 7481 6072
rect 7515 6069 7527 6103
rect 7469 6063 7527 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8352 6072 8861 6100
rect 8352 6060 8358 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 9646 6100 9674 6140
rect 10594 6128 10600 6140
rect 10652 6128 10658 6180
rect 10778 6100 10784 6112
rect 9646 6072 10784 6100
rect 8849 6063 8907 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11020 6072 11529 6100
rect 11020 6060 11026 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11624 6100 11652 6208
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13648 6236 13676 6264
rect 14384 6236 14412 6267
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 15764 6313 15792 6344
rect 16022 6332 16028 6344
rect 16080 6372 16086 6384
rect 17788 6381 17816 6412
rect 18156 6412 19800 6440
rect 17773 6375 17831 6381
rect 16080 6344 17448 6372
rect 16080 6332 16086 6344
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 14976 6276 15577 6304
rect 14976 6264 14982 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16129 6307 16187 6313
rect 16129 6273 16141 6307
rect 16175 6273 16187 6307
rect 16666 6304 16672 6316
rect 16579 6276 16672 6304
rect 16129 6267 16187 6273
rect 15470 6236 15476 6248
rect 13648 6208 14412 6236
rect 14936 6208 15476 6236
rect 14936 6180 14964 6208
rect 15470 6196 15476 6208
rect 15528 6236 15534 6248
rect 15856 6236 15884 6267
rect 15528 6208 15884 6236
rect 16132 6236 16160 6267
rect 16666 6264 16672 6276
rect 16724 6304 16730 6316
rect 17310 6304 17316 6316
rect 16724 6276 17316 6304
rect 16724 6264 16730 6276
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17420 6304 17448 6344
rect 17773 6341 17785 6375
rect 17819 6341 17831 6375
rect 17773 6335 17831 6341
rect 17954 6304 17960 6316
rect 17420 6276 17960 6304
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18156 6313 18184 6412
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 18230 6332 18236 6384
rect 18288 6372 18294 6384
rect 18288 6344 19012 6372
rect 18288 6332 18294 6344
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 18141 6267 18199 6273
rect 16574 6236 16580 6248
rect 16132 6208 16580 6236
rect 15528 6196 15534 6208
rect 16574 6196 16580 6208
rect 16632 6236 16638 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16632 6208 16773 6236
rect 16632 6196 16638 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 18064 6236 18092 6267
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18984 6313 19012 6344
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6273 19027 6307
rect 19518 6304 19524 6316
rect 19479 6276 19524 6304
rect 18969 6267 19027 6273
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 20530 6304 20536 6316
rect 20491 6276 20536 6304
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 18690 6236 18696 6248
rect 18064 6208 18696 6236
rect 16761 6199 16819 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 11974 6128 11980 6180
rect 12032 6168 12038 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12032 6140 12817 6168
rect 12032 6128 12038 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14458 6168 14464 6180
rect 14240 6140 14464 6168
rect 14240 6128 14246 6140
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 14918 6128 14924 6180
rect 14976 6128 14982 6180
rect 15933 6171 15991 6177
rect 15933 6137 15945 6171
rect 15979 6168 15991 6171
rect 20162 6168 20168 6180
rect 15979 6140 20168 6168
rect 15979 6137 15991 6140
rect 15933 6131 15991 6137
rect 20162 6128 20168 6140
rect 20220 6128 20226 6180
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11624 6072 11897 6100
rect 11517 6063 11575 6069
rect 11885 6069 11897 6072
rect 11931 6100 11943 6103
rect 12342 6100 12348 6112
rect 11931 6072 12348 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13722 6100 13728 6112
rect 13311 6072 13728 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 15010 6100 15016 6112
rect 14056 6072 15016 6100
rect 14056 6060 14062 6072
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 16025 6103 16083 6109
rect 16025 6100 16037 6103
rect 15252 6072 16037 6100
rect 15252 6060 15258 6072
rect 16025 6069 16037 6072
rect 16071 6100 16083 6103
rect 16298 6100 16304 6112
rect 16071 6072 16304 6100
rect 16071 6069 16083 6072
rect 16025 6063 16083 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 17126 6100 17132 6112
rect 16448 6072 17132 6100
rect 16448 6060 16454 6072
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 18414 6060 18420 6112
rect 18472 6100 18478 6112
rect 20070 6100 20076 6112
rect 18472 6072 20076 6100
rect 18472 6060 18478 6072
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20622 6100 20628 6112
rect 20583 6072 20628 6100
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 1104 6010 21436 6032
rect 1104 5958 4338 6010
rect 4390 5958 4402 6010
rect 4454 5958 4466 6010
rect 4518 5958 4530 6010
rect 4582 5958 4594 6010
rect 4646 5958 11116 6010
rect 11168 5958 11180 6010
rect 11232 5958 11244 6010
rect 11296 5958 11308 6010
rect 11360 5958 11372 6010
rect 11424 5958 17893 6010
rect 17945 5958 17957 6010
rect 18009 5958 18021 6010
rect 18073 5958 18085 6010
rect 18137 5958 18149 6010
rect 18201 5958 21436 6010
rect 1104 5936 21436 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2958 5896 2964 5908
rect 2919 5868 2964 5896
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 4982 5896 4988 5908
rect 4943 5868 4988 5896
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5316 5868 5917 5896
rect 5316 5856 5322 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 5905 5859 5963 5865
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7466 5896 7472 5908
rect 7423 5868 7472 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 16758 5896 16764 5908
rect 9364 5868 16764 5896
rect 9364 5856 9370 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 18414 5896 18420 5908
rect 17276 5868 18092 5896
rect 18375 5868 18420 5896
rect 17276 5856 17282 5868
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 2556 5800 3096 5828
rect 2556 5788 2562 5800
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 2958 5760 2964 5772
rect 2915 5732 2964 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 3068 5769 3096 5800
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 9582 5828 9588 5840
rect 5224 5800 6500 5828
rect 5224 5788 5230 5800
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5729 3111 5763
rect 5258 5760 5264 5772
rect 3053 5723 3111 5729
rect 4724 5732 5264 5760
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 3844 5664 4353 5692
rect 3844 5652 3850 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 4489 5695 4547 5701
rect 4489 5661 4501 5695
rect 4535 5692 4547 5695
rect 4724 5692 4752 5732
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 6472 5769 6500 5800
rect 9324 5800 9588 5828
rect 9324 5772 9352 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 18064 5828 18092 5868
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 18690 5896 18696 5908
rect 18651 5868 18696 5896
rect 18690 5856 18696 5868
rect 18748 5856 18754 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 19300 5868 19441 5896
rect 19300 5856 19306 5868
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 19978 5896 19984 5908
rect 19939 5868 19984 5896
rect 19429 5859 19487 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20622 5828 20628 5840
rect 9732 5800 18000 5828
rect 18064 5800 20628 5828
rect 9732 5788 9738 5800
rect 6457 5763 6515 5769
rect 5408 5732 6408 5760
rect 5408 5720 5414 5732
rect 4535 5664 4752 5692
rect 4535 5661 4547 5664
rect 4489 5655 4547 5661
rect 4798 5652 4804 5704
rect 4856 5701 4862 5704
rect 4856 5692 4864 5701
rect 6270 5692 6276 5704
rect 4856 5664 4901 5692
rect 6231 5664 6276 5692
rect 4856 5655 4864 5664
rect 4856 5652 4862 5655
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6380 5692 6408 5732
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 8021 5763 8079 5769
rect 6503 5732 7880 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 7466 5692 7472 5704
rect 6380 5664 7472 5692
rect 7466 5652 7472 5664
rect 7524 5692 7530 5704
rect 7650 5692 7656 5704
rect 7524 5664 7656 5692
rect 7524 5652 7530 5664
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7852 5692 7880 5732
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8570 5760 8576 5772
rect 8067 5732 8576 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9306 5720 9312 5772
rect 9364 5720 9370 5772
rect 9950 5760 9956 5772
rect 9416 5732 9956 5760
rect 9416 5701 9444 5732
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10652 5732 10793 5760
rect 10652 5720 10658 5732
rect 10781 5729 10793 5732
rect 10827 5760 10839 5763
rect 12710 5760 12716 5772
rect 10827 5732 12598 5760
rect 12671 5732 12716 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 9401 5695 9459 5701
rect 7852 5664 9260 5692
rect 2685 5627 2743 5633
rect 2685 5593 2697 5627
rect 2731 5624 2743 5627
rect 3694 5624 3700 5636
rect 2731 5596 3700 5624
rect 2731 5593 2743 5596
rect 2685 5587 2743 5593
rect 3694 5584 3700 5596
rect 3752 5584 3758 5636
rect 4617 5627 4675 5633
rect 4617 5593 4629 5627
rect 4663 5593 4675 5627
rect 4617 5587 4675 5593
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 3234 5556 3240 5568
rect 2823 5528 3240 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 4632 5556 4660 5587
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 4764 5596 4809 5624
rect 4764 5584 4770 5596
rect 4890 5584 4896 5636
rect 4948 5624 4954 5636
rect 7837 5627 7895 5633
rect 7837 5624 7849 5627
rect 4948 5596 7849 5624
rect 4948 5584 4954 5596
rect 7837 5593 7849 5596
rect 7883 5593 7895 5627
rect 9232 5624 9260 5664
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9582 5692 9588 5704
rect 9543 5664 9588 5692
rect 9401 5655 9459 5661
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 10410 5692 10416 5704
rect 9723 5664 10416 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 9232 5596 9444 5624
rect 7837 5587 7895 5593
rect 5350 5556 5356 5568
rect 4632 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6420 5528 6465 5556
rect 6420 5516 6426 5528
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7708 5528 7757 5556
rect 7708 5516 7714 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 9214 5556 9220 5568
rect 9175 5528 9220 5556
rect 7745 5519 7803 5525
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 9416 5556 9444 5596
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9692 5624 9720 5655
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10962 5692 10968 5704
rect 10551 5664 10968 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11112 5664 11529 5692
rect 11112 5652 11118 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11756 5664 11805 5692
rect 11756 5652 11762 5664
rect 11793 5661 11805 5664
rect 11839 5692 11851 5695
rect 11974 5692 11980 5704
rect 11839 5664 11980 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12570 5692 12598 5732
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13814 5760 13820 5772
rect 12943 5732 13820 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 12912 5692 12940 5723
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14424 5732 14565 5760
rect 14424 5720 14430 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 15010 5720 15016 5772
rect 15068 5760 15074 5772
rect 16485 5763 16543 5769
rect 16485 5760 16497 5763
rect 15068 5732 16497 5760
rect 15068 5720 15074 5732
rect 16485 5729 16497 5732
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 12570 5664 12940 5692
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 14090 5692 14096 5704
rect 13320 5664 14096 5692
rect 13320 5652 13326 5664
rect 14090 5652 14096 5664
rect 14148 5692 14154 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 14148 5664 14289 5692
rect 14148 5652 14154 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 14277 5655 14335 5661
rect 9548 5596 9720 5624
rect 9548 5584 9554 5596
rect 10686 5584 10692 5636
rect 10744 5624 10750 5636
rect 14292 5624 14320 5655
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 16022 5692 16028 5704
rect 15519 5664 16028 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16298 5702 16304 5704
rect 16224 5692 16304 5702
rect 16132 5664 16304 5692
rect 16132 5624 16160 5664
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 16574 5652 16580 5704
rect 16632 5692 16638 5704
rect 17586 5692 17592 5704
rect 16632 5664 16677 5692
rect 17547 5664 17592 5692
rect 16632 5652 16638 5664
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17972 5692 18000 5800
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5760 18475 5763
rect 18598 5760 18604 5772
rect 18463 5732 18604 5760
rect 18463 5729 18475 5732
rect 18417 5723 18475 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 20254 5720 20260 5772
rect 20312 5760 20318 5772
rect 20533 5763 20591 5769
rect 20533 5760 20545 5763
rect 20312 5732 20545 5760
rect 20312 5720 20318 5732
rect 20533 5729 20545 5732
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 18233 5695 18291 5701
rect 18233 5692 18245 5695
rect 17972 5664 18245 5692
rect 18233 5661 18245 5664
rect 18279 5661 18291 5695
rect 18506 5692 18512 5704
rect 18467 5664 18512 5692
rect 18233 5655 18291 5661
rect 10744 5596 11744 5624
rect 14292 5596 16160 5624
rect 18248 5624 18276 5655
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 19334 5692 19340 5704
rect 19295 5664 19340 5692
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20441 5695 20499 5701
rect 20441 5692 20453 5695
rect 20404 5664 20453 5692
rect 20404 5652 20410 5664
rect 20441 5661 20453 5664
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 18690 5624 18696 5636
rect 18248 5596 18696 5624
rect 10744 5584 10750 5596
rect 9950 5556 9956 5568
rect 9416 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 11716 5565 11744 5596
rect 18690 5584 18696 5596
rect 18748 5584 18754 5636
rect 10597 5559 10655 5565
rect 10597 5525 10609 5559
rect 10643 5556 10655 5559
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10643 5528 11345 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5525 11759 5559
rect 11701 5519 11759 5525
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12216 5528 12265 5556
rect 12216 5516 12222 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12253 5519 12311 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13688 5528 14105 5556
rect 13688 5516 13694 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 16117 5559 16175 5565
rect 16117 5525 16129 5559
rect 16163 5556 16175 5559
rect 17034 5556 17040 5568
rect 16163 5528 17040 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17681 5559 17739 5565
rect 17681 5525 17693 5559
rect 17727 5556 17739 5559
rect 18874 5556 18880 5568
rect 17727 5528 18880 5556
rect 17727 5525 17739 5528
rect 17681 5519 17739 5525
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 20162 5516 20168 5568
rect 20220 5556 20226 5568
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 20220 5528 20361 5556
rect 20220 5516 20226 5528
rect 20349 5525 20361 5528
rect 20395 5525 20407 5559
rect 20349 5519 20407 5525
rect 1104 5466 21436 5488
rect 1104 5414 7727 5466
rect 7779 5414 7791 5466
rect 7843 5414 7855 5466
rect 7907 5414 7919 5466
rect 7971 5414 7983 5466
rect 8035 5414 14504 5466
rect 14556 5414 14568 5466
rect 14620 5414 14632 5466
rect 14684 5414 14696 5466
rect 14748 5414 14760 5466
rect 14812 5414 21436 5466
rect 1104 5392 21436 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 3752 5324 5089 5352
rect 3752 5312 3758 5324
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6641 5355 6699 5361
rect 6641 5352 6653 5355
rect 6420 5324 6653 5352
rect 6420 5312 6426 5324
rect 6641 5321 6653 5324
rect 6687 5321 6699 5355
rect 6641 5315 6699 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9030 5352 9036 5364
rect 8987 5324 9036 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9272 5324 9965 5352
rect 9272 5312 9278 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 10781 5355 10839 5361
rect 10781 5321 10793 5355
rect 10827 5352 10839 5355
rect 11054 5352 11060 5364
rect 10827 5324 11060 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 1857 5287 1915 5293
rect 1857 5284 1869 5287
rect 1636 5256 1869 5284
rect 1636 5244 1642 5256
rect 1857 5253 1869 5256
rect 1903 5253 1915 5287
rect 7374 5284 7380 5296
rect 1857 5247 1915 5253
rect 6380 5256 7380 5284
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3050 5216 3056 5228
rect 3011 5188 3056 5216
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4154 5216 4160 5228
rect 4111 5188 4160 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5258 5216 5264 5228
rect 4939 5188 5264 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 4816 5148 4844 5179
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 6380 5225 6408 5256
rect 7374 5244 7380 5256
rect 7432 5284 7438 5296
rect 9674 5284 9680 5296
rect 7432 5256 7880 5284
rect 7432 5244 7438 5256
rect 6365 5219 6423 5225
rect 5408 5188 5453 5216
rect 5408 5176 5414 5188
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 6365 5179 6423 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7742 5216 7748 5228
rect 7607 5188 7748 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 7852 5225 7880 5256
rect 7944 5256 9680 5284
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 5368 5148 5396 5176
rect 4816 5120 5396 5148
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 6914 5148 6920 5160
rect 6687 5120 6920 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7944 5148 7972 5256
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 9858 5284 9864 5296
rect 9819 5256 9864 5284
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9122 5216 9128 5228
rect 8895 5188 9128 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9324 5216 9536 5222
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 9272 5194 10701 5216
rect 9272 5188 9352 5194
rect 9508 5188 10701 5194
rect 9272 5176 9278 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 9858 5148 9864 5160
rect 7024 5120 7972 5148
rect 9505 5140 9864 5148
rect 9324 5120 9864 5140
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 7024 5080 7052 5120
rect 9324 5112 9533 5120
rect 7650 5080 7656 5092
rect 4295 5052 7052 5080
rect 7611 5052 7656 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 9324 5080 9352 5112
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 9950 5108 9956 5160
rect 10008 5148 10014 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10008 5120 10149 5148
rect 10008 5108 10014 5120
rect 10137 5117 10149 5120
rect 10183 5148 10195 5151
rect 10594 5148 10600 5160
rect 10183 5120 10600 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 7892 5052 9352 5080
rect 7892 5040 7898 5052
rect 9582 5040 9588 5092
rect 9640 5080 9646 5092
rect 10796 5080 10824 5315
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 12618 5352 12624 5364
rect 12207 5324 12624 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13630 5352 13636 5364
rect 13591 5324 13636 5352
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 16669 5355 16727 5361
rect 13780 5324 13825 5352
rect 14292 5324 16528 5352
rect 13780 5312 13786 5324
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 11664 5256 11836 5284
rect 11664 5244 11670 5256
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11572 5188 11713 5216
rect 11572 5176 11578 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11808 5216 11836 5256
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 14292 5284 14320 5324
rect 12124 5256 14320 5284
rect 12124 5244 12130 5256
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 15933 5287 15991 5293
rect 14424 5256 15056 5284
rect 14424 5244 14430 5256
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 11808 5188 12357 5216
rect 11701 5179 11759 5185
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12584 5188 12633 5216
rect 12584 5176 12590 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 13964 5188 14473 5216
rect 13964 5176 13970 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 13446 5148 13452 5160
rect 11532 5120 13452 5148
rect 11532 5089 11560 5120
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13814 5148 13820 5160
rect 13775 5120 13820 5148
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14660 5148 14688 5179
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 14918 5216 14924 5228
rect 14792 5188 14924 5216
rect 14792 5176 14798 5188
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 15028 5225 15056 5256
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16206 5284 16212 5296
rect 15979 5256 16212 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 16500 5216 16528 5324
rect 16669 5321 16681 5355
rect 16715 5321 16727 5355
rect 17034 5352 17040 5364
rect 16995 5324 17040 5352
rect 16669 5315 16727 5321
rect 16684 5284 16712 5315
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 20346 5352 20352 5364
rect 18748 5324 19196 5352
rect 20307 5324 20352 5352
rect 18748 5312 18754 5324
rect 19058 5284 19064 5296
rect 16684 5256 19064 5284
rect 17678 5216 17684 5228
rect 16500 5188 17684 5216
rect 15013 5179 15071 5185
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 18892 5225 18920 5256
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5216 18107 5219
rect 18877 5219 18935 5225
rect 18095 5188 18828 5216
rect 18095 5185 18107 5188
rect 18049 5179 18107 5185
rect 14292 5120 14688 5148
rect 9640 5052 10824 5080
rect 11517 5083 11575 5089
rect 9640 5040 9646 5052
rect 11517 5049 11529 5083
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12529 5083 12587 5089
rect 12529 5080 12541 5083
rect 12400 5052 12541 5080
rect 12400 5040 12406 5052
rect 12529 5049 12541 5052
rect 12575 5080 12587 5083
rect 14182 5080 14188 5092
rect 12575 5052 14188 5080
rect 12575 5049 12587 5052
rect 12529 5043 12587 5049
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 6454 5012 6460 5024
rect 6415 4984 6460 5012
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7282 5012 7288 5024
rect 7064 4984 7288 5012
rect 7064 4972 7070 4984
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 9493 5015 9551 5021
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 9674 5012 9680 5024
rect 9539 4984 9680 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 13262 5012 13268 5024
rect 13223 4984 13268 5012
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 14292 5012 14320 5120
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 16264 5120 17141 5148
rect 16264 5108 16270 5120
rect 17129 5117 17141 5120
rect 17175 5117 17187 5151
rect 17129 5111 17187 5117
rect 17313 5151 17371 5157
rect 17313 5117 17325 5151
rect 17359 5148 17371 5151
rect 17494 5148 17500 5160
rect 17359 5120 17500 5148
rect 17359 5117 17371 5120
rect 17313 5111 17371 5117
rect 17494 5108 17500 5120
rect 17552 5108 17558 5160
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18380 5120 18705 5148
rect 18380 5108 18386 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18800 5148 18828 5188
rect 18877 5185 18889 5219
rect 18923 5185 18935 5219
rect 19168 5216 19196 5324
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 19245 5287 19303 5293
rect 19245 5253 19257 5287
rect 19291 5284 19303 5287
rect 19426 5284 19432 5296
rect 19291 5256 19432 5284
rect 19291 5253 19303 5256
rect 19245 5247 19303 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19889 5287 19947 5293
rect 19889 5253 19901 5287
rect 19935 5284 19947 5287
rect 20441 5287 20499 5293
rect 20441 5284 20453 5287
rect 19935 5256 20453 5284
rect 19935 5253 19947 5256
rect 19889 5247 19947 5253
rect 20088 5225 20116 5256
rect 20441 5253 20453 5256
rect 20487 5253 20499 5287
rect 20441 5247 20499 5253
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19168 5188 19993 5216
rect 18877 5179 18935 5185
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 20088 5219 20155 5225
rect 20088 5188 20109 5219
rect 19981 5179 20039 5185
rect 20097 5185 20109 5188
rect 20143 5185 20155 5219
rect 20097 5179 20155 5185
rect 19150 5148 19156 5160
rect 18800 5120 19156 5148
rect 18693 5111 18751 5117
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 19996 5148 20024 5179
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 19996 5120 20545 5148
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 17586 5080 17592 5092
rect 16163 5052 17592 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 17586 5040 17592 5052
rect 17644 5040 17650 5092
rect 18506 5040 18512 5092
rect 18564 5080 18570 5092
rect 18877 5083 18935 5089
rect 18877 5080 18889 5083
rect 18564 5052 18889 5080
rect 18564 5040 18570 5052
rect 18877 5049 18889 5052
rect 18923 5080 18935 5083
rect 19889 5083 19947 5089
rect 19889 5080 19901 5083
rect 18923 5052 19901 5080
rect 18923 5049 18935 5052
rect 18877 5043 18935 5049
rect 19889 5049 19901 5052
rect 19935 5049 19947 5083
rect 19889 5043 19947 5049
rect 13688 4984 14320 5012
rect 13688 4972 13694 4984
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14424 4984 14473 5012
rect 14424 4972 14430 4984
rect 14461 4981 14473 4984
rect 14507 4981 14519 5015
rect 14461 4975 14519 4981
rect 14921 5015 14979 5021
rect 14921 4981 14933 5015
rect 14967 5012 14979 5015
rect 15194 5012 15200 5024
rect 14967 4984 15200 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 21637 5015 21695 5021
rect 21637 5012 21649 5015
rect 18187 4984 21649 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 21637 4981 21649 4984
rect 21683 4981 21695 5015
rect 21637 4975 21695 4981
rect 1104 4922 21436 4944
rect 1104 4870 4338 4922
rect 4390 4870 4402 4922
rect 4454 4870 4466 4922
rect 4518 4870 4530 4922
rect 4582 4870 4594 4922
rect 4646 4870 11116 4922
rect 11168 4870 11180 4922
rect 11232 4870 11244 4922
rect 11296 4870 11308 4922
rect 11360 4870 11372 4922
rect 11424 4870 17893 4922
rect 17945 4870 17957 4922
rect 18009 4870 18021 4922
rect 18073 4870 18085 4922
rect 18137 4870 18149 4922
rect 18201 4870 21436 4922
rect 1104 4848 21436 4870
rect 3789 4811 3847 4817
rect 3789 4777 3801 4811
rect 3835 4808 3847 4811
rect 4890 4808 4896 4820
rect 3835 4780 4896 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6362 4808 6368 4820
rect 6227 4780 6368 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9398 4808 9404 4820
rect 9263 4780 9404 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 11333 4811 11391 4817
rect 11333 4808 11345 4811
rect 9640 4780 11345 4808
rect 9640 4768 9646 4780
rect 11333 4777 11345 4780
rect 11379 4777 11391 4811
rect 11333 4771 11391 4777
rect 15933 4811 15991 4817
rect 15933 4777 15945 4811
rect 15979 4808 15991 4811
rect 16206 4808 16212 4820
rect 15979 4780 16212 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 17037 4811 17095 4817
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17218 4808 17224 4820
rect 17083 4780 17224 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 18506 4768 18512 4820
rect 18564 4808 18570 4820
rect 18601 4811 18659 4817
rect 18601 4808 18613 4811
rect 18564 4780 18613 4808
rect 18564 4768 18570 4780
rect 18601 4777 18613 4780
rect 18647 4777 18659 4811
rect 18601 4771 18659 4777
rect 19794 4768 19800 4820
rect 19852 4808 19858 4820
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19852 4780 19901 4808
rect 19852 4768 19858 4780
rect 19889 4777 19901 4780
rect 19935 4777 19947 4811
rect 19889 4771 19947 4777
rect 5810 4740 5816 4752
rect 1688 4712 5816 4740
rect 1688 4681 1716 4712
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 9030 4700 9036 4752
rect 9088 4740 9094 4752
rect 9088 4712 10364 4740
rect 9088 4700 9094 4712
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4641 1731 4675
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 1673 4635 1731 4641
rect 4080 4644 4445 4672
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2682 4604 2688 4616
rect 1820 4576 2688 4604
rect 1820 4564 1826 4576
rect 2682 4564 2688 4576
rect 2740 4604 2746 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2740 4576 2881 4604
rect 2740 4564 2746 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3914 4607 3972 4613
rect 3914 4604 3926 4607
rect 3752 4576 3926 4604
rect 3752 4564 3758 4576
rect 3914 4573 3926 4576
rect 3960 4604 3972 4607
rect 4080 4604 4108 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9490 4672 9496 4684
rect 8987 4644 9496 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9490 4632 9496 4644
rect 9548 4672 9554 4684
rect 9953 4675 10011 4681
rect 9548 4644 9904 4672
rect 9548 4632 9554 4644
rect 3960 4576 4108 4604
rect 4341 4607 4399 4613
rect 3960 4573 3972 4576
rect 3914 4567 3972 4573
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 2590 4428 2596 4480
rect 2648 4468 2654 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 2648 4440 2697 4468
rect 2648 4428 2654 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 2685 4431 2743 4437
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3936 4440 3985 4468
rect 3936 4428 3942 4440
rect 3973 4437 3985 4440
rect 4019 4468 4031 4471
rect 4356 4468 4384 4567
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4764 4576 4905 4604
rect 4764 4564 4770 4576
rect 4893 4573 4905 4576
rect 4939 4604 4951 4607
rect 5350 4604 5356 4616
rect 4939 4576 5356 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5684 4576 6009 4604
rect 5684 4564 5690 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 5997 4567 6055 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6880 4576 7205 4604
rect 6880 4564 6886 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 9125 4607 9183 4613
rect 7800 4576 8984 4604
rect 7800 4564 7806 4576
rect 7006 4496 7012 4548
rect 7064 4536 7070 4548
rect 7834 4536 7840 4548
rect 7064 4508 7840 4536
rect 7064 4496 7070 4508
rect 7834 4496 7840 4508
rect 7892 4496 7898 4548
rect 8202 4536 8208 4548
rect 8163 4508 8208 4536
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 8846 4536 8852 4548
rect 8435 4508 8852 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 8956 4536 8984 4576
rect 9125 4573 9137 4607
rect 9171 4604 9183 4607
rect 9582 4604 9588 4616
rect 9171 4576 9588 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9876 4604 9904 4644
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10042 4672 10048 4684
rect 9999 4644 10048 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10152 4681 10180 4712
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10336 4672 10364 4712
rect 10502 4700 10508 4752
rect 10560 4740 10566 4752
rect 16945 4743 17003 4749
rect 16945 4740 16957 4743
rect 10560 4712 12940 4740
rect 10560 4700 10566 4712
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 10336 4644 11805 4672
rect 10137 4635 10195 4641
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12618 4672 12624 4684
rect 12207 4644 12624 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9876 4576 10241 4604
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10322 4607 10380 4613
rect 10322 4573 10334 4607
rect 10368 4573 10380 4607
rect 10322 4567 10380 4573
rect 8956 4508 9720 4536
rect 4019 4440 4384 4468
rect 4985 4471 5043 4477
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5074 4468 5080 4480
rect 5031 4440 5080 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 6365 4471 6423 4477
rect 6365 4437 6377 4471
rect 6411 4468 6423 4471
rect 6914 4468 6920 4480
rect 6411 4440 6920 4468
rect 6411 4437 6423 4440
rect 6365 4431 6423 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7285 4471 7343 4477
rect 7285 4468 7297 4471
rect 7156 4440 7297 4468
rect 7156 4428 7162 4440
rect 7285 4437 7297 4440
rect 7331 4437 7343 4471
rect 7285 4431 7343 4437
rect 9401 4471 9459 4477
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 9582 4468 9588 4480
rect 9447 4440 9588 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9692 4468 9720 4508
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 10336 4536 10364 4567
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 10965 4607 11023 4613
rect 10468 4576 10513 4604
rect 10468 4564 10474 4576
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11698 4604 11704 4616
rect 11011 4576 11704 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 9824 4508 10364 4536
rect 9824 4496 9830 4508
rect 10686 4496 10692 4548
rect 10744 4536 10750 4548
rect 11149 4539 11207 4545
rect 11149 4536 11161 4539
rect 10744 4508 11161 4536
rect 10744 4496 10750 4508
rect 11149 4505 11161 4508
rect 11195 4505 11207 4539
rect 11992 4536 12020 4567
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12250 4604 12256 4616
rect 12124 4576 12169 4604
rect 12211 4576 12256 4604
rect 12124 4564 12130 4576
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 12912 4613 12940 4712
rect 16132 4712 16957 4740
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 13044 4576 13093 4604
rect 13044 4564 13050 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 13412 4576 14565 4604
rect 13412 4564 13418 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 15194 4604 15200 4616
rect 14553 4567 14611 4573
rect 15120 4576 15200 4604
rect 12802 4536 12808 4548
rect 11992 4508 12808 4536
rect 11149 4499 11207 4505
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 15120 4536 15148 4576
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 16132 4613 16160 4712
rect 16945 4709 16957 4712
rect 16991 4740 17003 4743
rect 17589 4743 17647 4749
rect 17589 4740 17601 4743
rect 16991 4712 17601 4740
rect 16991 4709 17003 4712
rect 16945 4703 17003 4709
rect 17589 4709 17601 4712
rect 17635 4709 17647 4743
rect 17589 4703 17647 4709
rect 17678 4700 17684 4752
rect 17736 4740 17742 4752
rect 17736 4712 20576 4740
rect 17736 4700 17742 4712
rect 16482 4672 16488 4684
rect 16224 4644 16488 4672
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 12912 4508 15148 4536
rect 15289 4539 15347 4545
rect 12912 4468 12940 4508
rect 15289 4505 15301 4539
rect 15335 4536 15347 4539
rect 16224 4536 16252 4644
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 17402 4672 17408 4684
rect 17175 4644 17408 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 18656 4644 19288 4672
rect 18656 4632 18662 4644
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16666 4604 16672 4616
rect 16439 4576 16672 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 17862 4604 17868 4616
rect 17819 4576 17868 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 15335 4508 16252 4536
rect 16301 4539 16359 4545
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 16301 4505 16313 4539
rect 16347 4536 16359 4539
rect 16574 4536 16580 4548
rect 16347 4508 16580 4536
rect 16347 4505 16359 4508
rect 16301 4499 16359 4505
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16684 4536 16712 4564
rect 17604 4536 17632 4567
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18690 4604 18696 4616
rect 18651 4576 18696 4604
rect 18417 4567 18475 4573
rect 16684 4508 17632 4536
rect 18432 4536 18460 4567
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 19260 4613 19288 4644
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 20548 4613 20576 4712
rect 19710 4607 19768 4613
rect 19392 4576 19437 4604
rect 19392 4564 19398 4576
rect 19710 4573 19722 4607
rect 19756 4604 19768 4607
rect 20533 4607 20591 4613
rect 19756 4576 19840 4604
rect 19756 4573 19768 4576
rect 19710 4567 19768 4573
rect 19426 4536 19432 4548
rect 18432 4508 19432 4536
rect 19426 4496 19432 4508
rect 19484 4536 19490 4548
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 19484 4508 19533 4536
rect 19484 4496 19490 4508
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 19610 4496 19616 4548
rect 19668 4536 19674 4548
rect 19668 4508 19713 4536
rect 19668 4496 19674 4508
rect 9692 4440 12940 4468
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 13872 4440 14657 4468
rect 13872 4428 13878 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15381 4471 15439 4477
rect 15381 4468 15393 4471
rect 15252 4440 15393 4468
rect 15252 4428 15258 4440
rect 15381 4437 15393 4440
rect 15427 4437 15439 4471
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 15381 4431 15439 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 19150 4428 19156 4480
rect 19208 4468 19214 4480
rect 19812 4468 19840 4576
rect 20533 4573 20545 4607
rect 20579 4573 20591 4607
rect 20533 4567 20591 4573
rect 20714 4536 20720 4548
rect 20675 4508 20720 4536
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 19208 4440 19840 4468
rect 19208 4428 19214 4440
rect 1104 4378 21436 4400
rect 1104 4326 7727 4378
rect 7779 4326 7791 4378
rect 7843 4326 7855 4378
rect 7907 4326 7919 4378
rect 7971 4326 7983 4378
rect 8035 4326 14504 4378
rect 14556 4326 14568 4378
rect 14620 4326 14632 4378
rect 14684 4326 14696 4378
rect 14748 4326 14760 4378
rect 14812 4326 21436 4378
rect 1104 4304 21436 4326
rect 5534 4264 5540 4276
rect 1872 4236 5540 4264
rect 1872 4205 1900 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7282 4264 7288 4276
rect 7055 4236 7288 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 8573 4267 8631 4273
rect 8573 4233 8585 4267
rect 8619 4264 8631 4267
rect 9030 4264 9036 4276
rect 8619 4236 9036 4264
rect 8619 4233 8631 4236
rect 8573 4227 8631 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 15930 4264 15936 4276
rect 10928 4236 13768 4264
rect 15891 4236 15936 4264
rect 10928 4224 10934 4236
rect 1857 4199 1915 4205
rect 1857 4165 1869 4199
rect 1903 4165 1915 4199
rect 2590 4196 2596 4208
rect 2551 4168 2596 4196
rect 1857 4159 1915 4165
rect 2590 4156 2596 4168
rect 2648 4156 2654 4208
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 3752 4168 4016 4196
rect 3752 4156 3758 4168
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3988 4128 4016 4168
rect 5902 4156 5908 4208
rect 5960 4196 5966 4208
rect 5960 4168 6316 4196
rect 5960 4156 5966 4168
rect 4048 4131 4106 4137
rect 4048 4128 4060 4131
rect 3988 4100 4060 4128
rect 4048 4097 4060 4100
rect 4094 4097 4106 4131
rect 4048 4091 4106 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4433 4131 4491 4137
rect 4212 4100 4257 4128
rect 4212 4088 4218 4100
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4433 4091 4491 4097
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2866 4060 2872 4072
rect 2823 4032 2872 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4448 4060 4476 4091
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 6178 4128 6184 4140
rect 5675 4100 6184 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6288 4128 6316 4168
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 7745 4199 7803 4205
rect 6788 4168 7236 4196
rect 6788 4156 6794 4168
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6288 4100 6837 4128
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7208 4128 7236 4168
rect 7745 4165 7757 4199
rect 7791 4196 7803 4199
rect 8294 4196 8300 4208
rect 7791 4168 8300 4196
rect 7791 4165 7803 4168
rect 7745 4159 7803 4165
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 9692 4196 9720 4224
rect 10778 4196 10784 4208
rect 9692 4168 10088 4196
rect 10739 4168 10784 4196
rect 10060 4140 10088 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 12069 4199 12127 4205
rect 12069 4165 12081 4199
rect 12115 4196 12127 4199
rect 12894 4196 12900 4208
rect 12115 4168 12149 4196
rect 12855 4168 12900 4196
rect 12115 4165 12127 4168
rect 12069 4159 12127 4165
rect 8018 4128 8024 4140
rect 7208 4100 8024 4128
rect 7101 4091 7159 4097
rect 5074 4060 5080 4072
rect 4304 4032 5080 4060
rect 4304 4020 4310 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 5132 4032 6653 4060
rect 5132 4020 5138 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 3329 3995 3387 4001
rect 2087 3964 2774 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 2746 3936 2774 3964
rect 3329 3961 3341 3995
rect 3375 3992 3387 3995
rect 3970 3992 3976 4004
rect 3375 3964 3976 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 3970 3952 3976 3964
rect 4028 3992 4034 4004
rect 4341 3995 4399 4001
rect 4341 3992 4353 3995
rect 4028 3964 4353 3992
rect 4028 3952 4034 3964
rect 4341 3961 4353 3964
rect 4387 3961 4399 3995
rect 4341 3955 4399 3961
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5442 3992 5448 4004
rect 4764 3964 5448 3992
rect 4764 3952 4770 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5721 3995 5779 4001
rect 5721 3961 5733 3995
rect 5767 3992 5779 3995
rect 7116 3992 7144 4091
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8570 4131 8628 4137
rect 8570 4097 8582 4131
rect 8616 4128 8628 4131
rect 9674 4131 9732 4137
rect 8616 4100 9076 4128
rect 8616 4097 8628 4100
rect 8570 4091 8628 4097
rect 9048 4069 9076 4100
rect 9674 4097 9686 4131
rect 9720 4128 9732 4131
rect 10042 4128 10048 4140
rect 9720 4100 9904 4128
rect 9955 4100 10048 4128
rect 9720 4097 9732 4100
rect 9674 4091 9732 4097
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4060 9091 4063
rect 9766 4060 9772 4072
rect 9079 4032 9772 4060
rect 9079 4029 9091 4032
rect 9033 4023 9091 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9876 4060 9904 4100
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10318 4128 10324 4140
rect 10183 4100 10324 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10152 4060 10180 4091
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12084 4128 12112 4159
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 13740 4205 13768 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17037 4267 17095 4273
rect 16632 4236 16988 4264
rect 16632 4224 16638 4236
rect 13725 4199 13783 4205
rect 13725 4165 13737 4199
rect 13771 4165 13783 4199
rect 16850 4196 16856 4208
rect 13725 4159 13783 4165
rect 16040 4168 16856 4196
rect 12618 4128 12624 4140
rect 11839 4100 12434 4128
rect 12579 4100 12624 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 9876 4032 10180 4060
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 11698 4060 11704 4072
rect 11655 4032 11704 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 11698 4020 11704 4032
rect 11756 4060 11762 4072
rect 12066 4060 12072 4072
rect 11756 4032 12072 4060
rect 11756 4020 11762 4032
rect 12066 4020 12072 4032
rect 12124 4060 12130 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 12124 4032 12173 4060
rect 12124 4020 12130 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 7282 3992 7288 4004
rect 5767 3964 7288 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 9398 3992 9404 4004
rect 7975 3964 9404 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 10612 3964 11468 3992
rect 2746 3896 2780 3936
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4120 3896 5089 3924
rect 4120 3884 4126 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 5077 3887 5135 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 6696 3896 6745 3924
rect 6696 3884 6702 3896
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8352 3896 8401 3924
rect 8352 3884 8358 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8941 3927 8999 3933
rect 8941 3893 8953 3927
rect 8987 3924 8999 3927
rect 9030 3924 9036 3936
rect 8987 3896 9036 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 10612 3924 10640 3964
rect 9180 3896 10640 3924
rect 9180 3884 9186 3896
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 10873 3927 10931 3933
rect 10873 3924 10885 3927
rect 10744 3896 10885 3924
rect 10744 3884 10750 3896
rect 10873 3893 10885 3896
rect 10919 3893 10931 3927
rect 11440 3924 11468 3964
rect 11514 3952 11520 4004
rect 11572 3992 11578 4004
rect 12406 3992 12434 4100
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12802 4128 12808 4140
rect 12715 4100 12808 4128
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13262 4128 13268 4140
rect 13035 4100 13268 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 13504 4100 14657 4128
rect 13504 4088 13510 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 15102 4088 15108 4140
rect 15160 4128 15166 4140
rect 15657 4131 15715 4137
rect 15657 4128 15669 4131
rect 15160 4100 15669 4128
rect 15160 4088 15166 4100
rect 15657 4097 15669 4100
rect 15703 4097 15715 4131
rect 15657 4091 15715 4097
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4128 15807 4131
rect 15838 4128 15844 4140
rect 15795 4100 15844 4128
rect 15795 4097 15807 4100
rect 15749 4091 15807 4097
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16040 4137 16068 4168
rect 16850 4156 16856 4168
rect 16908 4156 16914 4208
rect 16960 4196 16988 4236
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 17402 4264 17408 4276
rect 17083 4236 17408 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 19150 4264 19156 4276
rect 17972 4236 19156 4264
rect 17862 4196 17868 4208
rect 16960 4168 17868 4196
rect 16025 4131 16083 4137
rect 16025 4128 16037 4131
rect 15988 4100 16037 4128
rect 15988 4088 15994 4100
rect 16025 4097 16037 4100
rect 16071 4097 16083 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 16025 4091 16083 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4128 16819 4131
rect 16960 4128 16988 4168
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 17972 4205 18000 4236
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 17957 4199 18015 4205
rect 17957 4165 17969 4199
rect 18003 4165 18015 4199
rect 17957 4159 18015 4165
rect 18141 4199 18199 4205
rect 18141 4165 18153 4199
rect 18187 4196 18199 4199
rect 19061 4199 19119 4205
rect 19061 4196 19073 4199
rect 18187 4168 19073 4196
rect 18187 4165 18199 4168
rect 18141 4159 18199 4165
rect 19061 4165 19073 4168
rect 19107 4196 19119 4199
rect 19610 4196 19616 4208
rect 19107 4168 19616 4196
rect 19107 4165 19119 4168
rect 19061 4159 19119 4165
rect 16807 4100 16988 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 12820 4060 12848 4088
rect 14734 4060 14740 4072
rect 12820 4032 14740 4060
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 16574 4060 16580 4072
rect 14875 4032 16580 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 13173 3995 13231 4001
rect 13173 3992 13185 3995
rect 11572 3964 12020 3992
rect 12406 3964 13185 3992
rect 11572 3952 11578 3964
rect 11606 3924 11612 3936
rect 11440 3896 11612 3924
rect 10873 3887 10931 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11848 3896 11897 3924
rect 11848 3884 11854 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11992 3924 12020 3964
rect 13173 3961 13185 3964
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 18156 3992 18184 4159
rect 19610 4156 19616 4168
rect 19668 4196 19674 4208
rect 19889 4199 19947 4205
rect 19889 4196 19901 4199
rect 19668 4168 19901 4196
rect 19668 4156 19674 4168
rect 19889 4165 19901 4168
rect 19935 4165 19947 4199
rect 19889 4159 19947 4165
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18288 4100 18797 4128
rect 18288 4088 18294 4100
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4097 19027 4131
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 18969 4091 19027 4097
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 18984 4060 19012 4091
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19702 4088 19708 4140
rect 19760 4128 19766 4140
rect 19797 4131 19855 4137
rect 19797 4128 19809 4131
rect 19760 4100 19809 4128
rect 19760 4088 19766 4100
rect 19797 4097 19809 4100
rect 19843 4097 19855 4131
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 19797 4091 19855 4097
rect 20254 4088 20260 4100
rect 20312 4128 20318 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20312 4100 20545 4128
rect 20312 4088 20318 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 20533 4091 20591 4097
rect 19334 4060 19340 4072
rect 18371 4032 19340 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 15611 3964 18184 3992
rect 20717 3995 20775 4001
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 20717 3961 20729 3995
rect 20763 3992 20775 3995
rect 20806 3992 20812 4004
rect 20763 3964 20812 3992
rect 20763 3961 20775 3964
rect 20717 3955 20775 3961
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 12986 3924 12992 3936
rect 11992 3896 12992 3924
rect 11885 3887 11943 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13136 3896 13829 3924
rect 13136 3884 13142 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15252 3896 15301 3924
rect 15252 3884 15258 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 16758 3924 16764 3936
rect 16719 3896 16764 3924
rect 15289 3887 15347 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 19337 3927 19395 3933
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 20070 3924 20076 3936
rect 19383 3896 20076 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21637 3927 21695 3933
rect 21637 3924 21649 3927
rect 21416 3896 21649 3924
rect 21416 3884 21422 3896
rect 21637 3893 21649 3896
rect 21683 3893 21695 3927
rect 21637 3887 21695 3893
rect 1104 3834 21436 3856
rect 1104 3782 4338 3834
rect 4390 3782 4402 3834
rect 4454 3782 4466 3834
rect 4518 3782 4530 3834
rect 4582 3782 4594 3834
rect 4646 3782 11116 3834
rect 11168 3782 11180 3834
rect 11232 3782 11244 3834
rect 11296 3782 11308 3834
rect 11360 3782 11372 3834
rect 11424 3782 17893 3834
rect 17945 3782 17957 3834
rect 18009 3782 18021 3834
rect 18073 3782 18085 3834
rect 18137 3782 18149 3834
rect 18201 3782 21436 3834
rect 1104 3760 21436 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3694 3720 3700 3732
rect 3016 3692 3700 3720
rect 3016 3680 3022 3692
rect 3694 3680 3700 3692
rect 3752 3720 3758 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 3752 3692 4445 3720
rect 3752 3680 3758 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 5592 3692 6101 3720
rect 5592 3680 5598 3692
rect 6089 3689 6101 3692
rect 6135 3720 6147 3723
rect 6454 3720 6460 3732
rect 6135 3692 6460 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7650 3720 7656 3732
rect 7239 3692 7656 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9766 3720 9772 3732
rect 9355 3692 9772 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10134 3720 10140 3732
rect 9907 3692 10140 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10410 3720 10416 3732
rect 10371 3692 10416 3720
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 11698 3720 11704 3732
rect 11659 3692 11704 3720
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 12216 3692 12265 3720
rect 12216 3680 12222 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12676 3692 12909 3720
rect 12676 3680 12682 3692
rect 12897 3689 12909 3692
rect 12943 3720 12955 3723
rect 14274 3720 14280 3732
rect 12943 3692 14280 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 14274 3680 14280 3692
rect 14332 3720 14338 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14332 3692 14657 3720
rect 14332 3680 14338 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15344 3692 15669 3720
rect 15344 3680 15350 3692
rect 15657 3689 15669 3692
rect 15703 3689 15715 3723
rect 15657 3683 15715 3689
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17770 3720 17776 3732
rect 16632 3692 17776 3720
rect 16632 3680 16638 3692
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18414 3720 18420 3732
rect 18375 3692 18420 3720
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 4246 3652 4252 3664
rect 4080 3624 4252 3652
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 3970 3516 3976 3528
rect 3927 3488 3976 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4080 3525 4108 3624
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 5350 3652 5356 3664
rect 4396 3624 5356 3652
rect 4396 3612 4402 3624
rect 5350 3612 5356 3624
rect 5408 3652 5414 3664
rect 5408 3624 6868 3652
rect 5408 3612 5414 3624
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5224 3556 5457 3584
rect 5224 3544 5230 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5718 3584 5724 3596
rect 5445 3547 5503 3553
rect 5552 3556 5724 3584
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4522 3516 4528 3528
rect 4295 3488 4528 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5552 3516 5580 3556
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5000 3488 5580 3516
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 1544 3420 1869 3448
rect 1544 3408 1550 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 3050 3448 3056 3460
rect 3011 3420 3056 3448
rect 1857 3411 1915 3417
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 4154 3448 4160 3460
rect 4067 3420 4160 3448
rect 4154 3408 4160 3420
rect 4212 3448 4218 3460
rect 4338 3448 4344 3460
rect 4212 3420 4344 3448
rect 4212 3408 4218 3420
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 5000 3448 5028 3488
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5684 3488 6101 3516
rect 5684 3476 5690 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 6236 3488 6285 3516
rect 6236 3476 6242 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6420 3488 6745 3516
rect 6420 3476 6426 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6840 3516 6868 3624
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 6972 3624 13216 3652
rect 6972 3612 6978 3624
rect 8205 3587 8263 3593
rect 8205 3584 8217 3587
rect 7300 3556 8217 3584
rect 7300 3528 7328 3556
rect 8205 3553 8217 3556
rect 8251 3553 8263 3587
rect 9674 3584 9680 3596
rect 8205 3547 8263 3553
rect 8404 3556 9680 3584
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6840 3488 6929 3516
rect 6733 3479 6791 3485
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7282 3516 7288 3528
rect 7064 3488 7109 3516
rect 7243 3488 7288 3516
rect 7064 3476 7070 3488
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7432 3488 7941 3516
rect 7432 3476 7438 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 8076 3488 8125 3516
rect 8076 3476 8082 3488
rect 8113 3485 8125 3488
rect 8159 3516 8171 3519
rect 8404 3516 8432 3556
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10100 3556 11069 3584
rect 10100 3544 10106 3556
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 12066 3584 12072 3596
rect 11057 3547 11115 3553
rect 11897 3556 12072 3584
rect 8159 3488 8432 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9490 3519 9548 3525
rect 9490 3516 9502 3519
rect 9364 3488 9502 3516
rect 9364 3476 9370 3488
rect 9490 3485 9502 3488
rect 9536 3516 9548 3519
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9536 3488 9965 3516
rect 9536 3485 9548 3488
rect 9490 3479 9548 3485
rect 9953 3485 9965 3488
rect 9999 3516 10011 3519
rect 10226 3516 10232 3528
rect 9999 3488 10232 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10502 3476 10508 3528
rect 10560 3516 10566 3528
rect 11897 3525 11925 3556
rect 12066 3544 12072 3556
rect 12124 3584 12130 3596
rect 12342 3584 12348 3596
rect 12124 3556 12348 3584
rect 12124 3544 12130 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 13188 3584 13216 3624
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13449 3655 13507 3661
rect 13449 3652 13461 3655
rect 13320 3624 13461 3652
rect 13320 3612 13326 3624
rect 13449 3621 13461 3624
rect 13495 3621 13507 3655
rect 13449 3615 13507 3621
rect 13906 3612 13912 3664
rect 13964 3652 13970 3664
rect 15010 3652 15016 3664
rect 13964 3624 15016 3652
rect 13964 3612 13970 3624
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 16666 3652 16672 3664
rect 15580 3624 16672 3652
rect 15580 3584 15608 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 17037 3655 17095 3661
rect 17037 3621 17049 3655
rect 17083 3652 17095 3655
rect 18325 3655 18383 3661
rect 18325 3652 18337 3655
rect 17083 3624 18337 3652
rect 17083 3621 17095 3624
rect 17037 3615 17095 3621
rect 18325 3621 18337 3624
rect 18371 3652 18383 3655
rect 18598 3652 18604 3664
rect 18371 3624 18604 3652
rect 18371 3621 18383 3624
rect 18325 3615 18383 3621
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 20717 3655 20775 3661
rect 20717 3621 20729 3655
rect 20763 3652 20775 3655
rect 21545 3655 21603 3661
rect 21545 3652 21557 3655
rect 20763 3624 21557 3652
rect 20763 3621 20775 3624
rect 20717 3615 20775 3621
rect 21545 3621 21557 3624
rect 21591 3621 21603 3655
rect 21545 3615 21603 3621
rect 13188 3556 15608 3584
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17276 3556 17509 3584
rect 17276 3544 17282 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17497 3547 17555 3553
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3584 17739 3587
rect 17862 3584 17868 3596
rect 17727 3556 17868 3584
rect 17727 3553 17739 3556
rect 17681 3547 17739 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 19334 3584 19340 3596
rect 18555 3556 19340 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10560 3488 10609 3516
rect 10560 3476 10566 3488
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 11882 3519 11940 3525
rect 10735 3488 11100 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 4448 3420 5028 3448
rect 5261 3451 5319 3457
rect 14 3340 20 3392
rect 72 3380 78 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 72 3352 1961 3380
rect 72 3340 78 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 1949 3343 2007 3349
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 3145 3383 3203 3389
rect 3145 3380 3157 3383
rect 2280 3352 3157 3380
rect 2280 3340 2286 3352
rect 3145 3349 3157 3352
rect 3191 3349 3203 3383
rect 3145 3343 3203 3349
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4448 3380 4476 3420
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 5307 3420 7757 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 10244 3448 10272 3476
rect 10781 3451 10839 3457
rect 10781 3448 10793 3451
rect 10244 3420 10793 3448
rect 7745 3411 7803 3417
rect 10781 3417 10793 3420
rect 10827 3417 10839 3451
rect 10781 3411 10839 3417
rect 10870 3408 10876 3460
rect 10928 3457 10934 3460
rect 10928 3451 10957 3457
rect 10945 3417 10957 3451
rect 10928 3411 10957 3417
rect 10928 3408 10934 3411
rect 4028 3352 4476 3380
rect 4028 3340 4034 3352
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 4798 3380 4804 3392
rect 4580 3352 4804 3380
rect 4580 3340 4586 3352
rect 4798 3340 4804 3352
rect 4856 3380 4862 3392
rect 4893 3383 4951 3389
rect 4893 3380 4905 3383
rect 4856 3352 4905 3380
rect 4856 3340 4862 3352
rect 4893 3349 4905 3352
rect 4939 3349 4951 3383
rect 4893 3343 4951 3349
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 6733 3383 6791 3389
rect 5408 3352 5453 3380
rect 5408 3340 5414 3352
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7006 3380 7012 3392
rect 6779 3352 7012 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 9674 3380 9680 3392
rect 9539 3352 9680 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 9674 3340 9680 3352
rect 9732 3380 9738 3392
rect 10134 3380 10140 3392
rect 9732 3352 10140 3380
rect 9732 3340 9738 3352
rect 10134 3340 10140 3352
rect 10192 3380 10198 3392
rect 11072 3380 11100 3488
rect 11882 3485 11894 3519
rect 11928 3485 11940 3519
rect 11882 3479 11940 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12032 3488 12817 3516
rect 12032 3476 12038 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 13078 3519 13136 3525
rect 13078 3516 13090 3519
rect 12952 3488 13090 3516
rect 12952 3476 12958 3488
rect 13078 3485 13090 3488
rect 13124 3516 13136 3519
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13124 3488 13553 3516
rect 13124 3485 13136 3488
rect 13078 3479 13136 3485
rect 13541 3485 13553 3488
rect 13587 3516 13599 3519
rect 13630 3516 13636 3528
rect 13587 3488 13636 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14274 3519 14332 3525
rect 14274 3485 14286 3519
rect 14320 3516 14332 3519
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14320 3488 14749 3516
rect 14320 3485 14332 3488
rect 14274 3479 14332 3485
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 14826 3516 14832 3528
rect 14783 3488 14832 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15194 3516 15200 3528
rect 15155 3488 15200 3516
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15749 3519 15807 3525
rect 15528 3488 15573 3516
rect 15528 3476 15534 3488
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 15930 3516 15936 3528
rect 15795 3488 15936 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 17954 3516 17960 3528
rect 16224 3488 17960 3516
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 16224 3448 16252 3488
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 18196 3488 18245 3516
rect 18196 3476 18202 3488
rect 18233 3485 18245 3488
rect 18279 3516 18291 3519
rect 19702 3516 19708 3528
rect 18279 3488 19708 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 16390 3448 16396 3460
rect 11664 3420 16252 3448
rect 16351 3420 16396 3448
rect 11664 3408 11670 3420
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 16577 3451 16635 3457
rect 16577 3417 16589 3451
rect 16623 3448 16635 3451
rect 19518 3448 19524 3460
rect 16623 3420 18368 3448
rect 19479 3420 19524 3448
rect 16623 3417 16635 3420
rect 16577 3411 16635 3417
rect 18340 3392 18368 3420
rect 19518 3408 19524 3420
rect 19576 3448 19582 3460
rect 19797 3451 19855 3457
rect 19797 3448 19809 3451
rect 19576 3420 19809 3448
rect 19576 3408 19582 3420
rect 19797 3417 19809 3420
rect 19843 3417 19855 3451
rect 19978 3448 19984 3460
rect 19939 3420 19984 3448
rect 19797 3411 19855 3417
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 20533 3451 20591 3457
rect 20533 3417 20545 3451
rect 20579 3448 20591 3451
rect 21910 3448 21916 3460
rect 20579 3420 21916 3448
rect 20579 3417 20591 3420
rect 20533 3411 20591 3417
rect 21910 3408 21916 3420
rect 21968 3408 21974 3460
rect 10192 3352 11100 3380
rect 11885 3383 11943 3389
rect 10192 3340 10198 3352
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 12158 3380 12164 3392
rect 11931 3352 12164 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 12851 3352 13093 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 13081 3349 13093 3352
rect 13127 3380 13139 3383
rect 13262 3380 13268 3392
rect 13127 3352 13268 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 15654 3380 15660 3392
rect 15243 3352 15660 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 17402 3380 17408 3392
rect 17363 3352 17408 3380
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 17862 3380 17868 3392
rect 17552 3352 17868 3380
rect 17552 3340 17558 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 18322 3340 18328 3392
rect 18380 3340 18386 3392
rect 1104 3290 21436 3312
rect 1104 3238 7727 3290
rect 7779 3238 7791 3290
rect 7843 3238 7855 3290
rect 7907 3238 7919 3290
rect 7971 3238 7983 3290
rect 8035 3238 14504 3290
rect 14556 3238 14568 3290
rect 14620 3238 14632 3290
rect 14684 3238 14696 3290
rect 14748 3238 14760 3290
rect 14812 3238 21436 3290
rect 1104 3216 21436 3238
rect 1486 3176 1492 3188
rect 1447 3148 1492 3176
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 5261 3179 5319 3185
rect 4111 3148 5212 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 2130 3068 2136 3120
rect 2188 3108 2194 3120
rect 2225 3111 2283 3117
rect 2225 3108 2237 3111
rect 2188 3080 2237 3108
rect 2188 3068 2194 3080
rect 2225 3077 2237 3080
rect 2271 3077 2283 3111
rect 2225 3071 2283 3077
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 3142 3108 3148 3120
rect 3099 3080 3148 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 3786 3068 3792 3120
rect 3844 3108 3850 3120
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 3844 3080 4169 3108
rect 3844 3068 3850 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2682 3040 2688 3052
rect 1719 3012 2688 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3694 3040 3700 3052
rect 3655 3012 3700 3040
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3896 3049 3924 3080
rect 4157 3077 4169 3080
rect 4203 3077 4215 3111
rect 5184 3108 5212 3148
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5350 3176 5356 3188
rect 5307 3148 5356 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6178 3176 6184 3188
rect 5675 3148 6184 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 9582 3176 9588 3188
rect 8444 3148 8892 3176
rect 9543 3148 9588 3176
rect 8444 3136 8450 3148
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 5184 3080 7113 3108
rect 4157 3071 4215 3077
rect 7101 3077 7113 3080
rect 7147 3077 7159 3111
rect 7101 3071 7159 3077
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 7340 3080 8432 3108
rect 7340 3068 7346 3080
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 5445 3043 5503 3049
rect 3927 3012 3961 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 5445 3009 5457 3043
rect 5491 3040 5503 3043
rect 5534 3040 5540 3052
rect 5491 3012 5540 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5684 3012 5733 3040
rect 5684 3000 5690 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 8205 3043 8263 3049
rect 5721 3003 5779 3009
rect 7116 3012 8156 3040
rect 3712 2972 3740 3000
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 2746 2944 3648 2972
rect 3712 2944 4261 2972
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 624 2876 2452 2904
rect 624 2864 630 2876
rect 1118 2796 1124 2848
rect 1176 2836 1182 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1176 2808 2329 2836
rect 1176 2796 1182 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2424 2836 2452 2876
rect 2746 2836 2774 2944
rect 3237 2907 3295 2913
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 3510 2904 3516 2916
rect 3283 2876 3516 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 3620 2904 3648 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4890 2972 4896 2984
rect 4249 2935 4307 2941
rect 4356 2944 4896 2972
rect 4356 2904 4384 2944
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 7116 2972 7144 3012
rect 7282 2972 7288 2984
rect 5040 2944 7144 2972
rect 7243 2944 7288 2972
rect 5040 2932 5046 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 8128 2972 8156 3012
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 8294 3040 8300 3052
rect 8251 3012 8300 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8404 2981 8432 3080
rect 8389 2975 8447 2981
rect 8128 2944 8340 2972
rect 3620 2876 4384 2904
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 8202 2904 8208 2916
rect 6687 2876 8208 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 2424 2808 2774 2836
rect 2317 2799 2375 2805
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 3108 2808 7849 2836
rect 3108 2796 3114 2808
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 8312 2836 8340 2944
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 8570 2972 8576 2984
rect 8435 2944 8576 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 8864 2972 8892 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10502 3176 10508 3188
rect 10463 3148 10508 3176
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 12069 3179 12127 3185
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 12250 3176 12256 3188
rect 12115 3148 12256 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12434 3136 12440 3188
rect 12492 3136 12498 3188
rect 12526 3136 12532 3188
rect 12584 3142 12590 3188
rect 12584 3136 12598 3142
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14148 3148 14565 3176
rect 14148 3136 14154 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 14553 3139 14611 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 15749 3179 15807 3185
rect 15749 3145 15761 3179
rect 15795 3176 15807 3179
rect 17957 3179 18015 3185
rect 17957 3176 17969 3179
rect 15795 3148 17969 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 17957 3145 17969 3148
rect 18003 3145 18015 3179
rect 17957 3139 18015 3145
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 18230 3176 18236 3188
rect 18187 3148 18236 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 9217 3111 9275 3117
rect 9217 3077 9229 3111
rect 9263 3108 9275 3111
rect 9766 3108 9772 3120
rect 9263 3080 9772 3108
rect 9263 3077 9275 3080
rect 9217 3071 9275 3077
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 10137 3111 10195 3117
rect 10137 3108 10149 3111
rect 10100 3080 10149 3108
rect 10100 3068 10106 3080
rect 10137 3077 10149 3080
rect 10183 3077 10195 3111
rect 10318 3108 10324 3120
rect 10279 3080 10324 3108
rect 10137 3071 10195 3077
rect 10318 3068 10324 3080
rect 10376 3108 10382 3120
rect 10870 3108 10876 3120
rect 10376 3080 10876 3108
rect 10376 3068 10382 3080
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 11974 3068 11980 3120
rect 12032 3108 12038 3120
rect 12346 3111 12404 3117
rect 12346 3108 12358 3111
rect 12032 3080 12358 3108
rect 12032 3068 12038 3080
rect 12346 3077 12358 3080
rect 12392 3077 12404 3111
rect 12346 3071 12404 3077
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 9674 3040 9680 3052
rect 9447 3012 9680 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 12452 3049 12480 3136
rect 12544 3117 12598 3136
rect 12544 3114 12613 3117
rect 12555 3111 12613 3114
rect 12555 3077 12567 3111
rect 12601 3077 12613 3111
rect 12555 3071 12613 3077
rect 12802 3068 12808 3120
rect 12860 3108 12866 3120
rect 13541 3111 13599 3117
rect 13541 3108 13553 3111
rect 12860 3080 13553 3108
rect 12860 3068 12866 3080
rect 13541 3077 13553 3080
rect 13587 3077 13599 3111
rect 13541 3071 13599 3077
rect 14366 3068 14372 3120
rect 14424 3108 14430 3120
rect 14461 3111 14519 3117
rect 14461 3108 14473 3111
rect 14424 3080 14473 3108
rect 14424 3068 14430 3080
rect 14461 3077 14473 3080
rect 14507 3077 14519 3111
rect 16485 3111 16543 3117
rect 16485 3108 16497 3111
rect 14461 3071 14519 3077
rect 14568 3080 16497 3108
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3009 12495 3043
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 12437 3003 12495 3009
rect 9858 2972 9864 2984
rect 8864 2944 9864 2972
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 12268 2972 12296 3003
rect 12710 3000 12716 3012
rect 12768 3040 12774 3052
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 12768 3012 13185 3040
rect 12768 3000 12774 3012
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13354 3040 13360 3052
rect 13315 3012 13360 3040
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 14568 3040 14596 3080
rect 16485 3077 16497 3080
rect 16531 3077 16543 3111
rect 16485 3071 16543 3077
rect 16761 3111 16819 3117
rect 16761 3077 16773 3111
rect 16807 3108 16819 3111
rect 17402 3108 17408 3120
rect 16807 3080 17408 3108
rect 16807 3077 16819 3080
rect 16761 3071 16819 3077
rect 17402 3068 17408 3080
rect 17460 3068 17466 3120
rect 20625 3111 20683 3117
rect 20625 3108 20637 3111
rect 17512 3080 20637 3108
rect 13688 3012 14596 3040
rect 13688 3000 13694 3012
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 15068 3012 16681 3040
rect 15068 3000 15074 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 16669 3003 16727 3009
rect 16776 3012 16957 3040
rect 14737 2975 14795 2981
rect 12268 2944 12388 2972
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 12158 2904 12164 2916
rect 8812 2876 12164 2904
rect 8812 2864 8818 2876
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12360 2904 12388 2944
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 14783 2944 15853 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15841 2941 15853 2944
rect 15887 2972 15899 2975
rect 16114 2972 16120 2984
rect 15887 2944 16120 2972
rect 15887 2941 15899 2944
rect 15841 2935 15899 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 16776 2972 16804 3012
rect 16945 3009 16957 3012
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17512 3040 17540 3080
rect 20625 3077 20637 3080
rect 20671 3077 20683 3111
rect 20625 3071 20683 3077
rect 17184 3012 17540 3040
rect 18138 3043 18196 3049
rect 17184 3000 17190 3012
rect 18138 3009 18150 3043
rect 18184 3009 18196 3043
rect 18138 3003 18196 3009
rect 16356 2944 16804 2972
rect 16356 2932 16362 2944
rect 16850 2932 16856 2984
rect 16908 2972 16914 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16908 2944 17233 2972
rect 16908 2932 16914 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 18156 2972 18184 3003
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18288 3012 18521 3040
rect 18288 3000 18294 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 19702 3040 19708 3052
rect 19663 3012 19708 3040
rect 18509 3003 18567 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20312 3012 20453 3040
rect 20312 3000 20318 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 18414 2972 18420 2984
rect 18156 2944 18420 2972
rect 17221 2935 17279 2941
rect 18414 2932 18420 2944
rect 18472 2972 18478 2984
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 18472 2944 18613 2972
rect 18472 2932 18478 2944
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 18601 2935 18659 2941
rect 12434 2904 12440 2916
rect 12360 2876 12440 2904
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 15289 2907 15347 2913
rect 15289 2904 15301 2907
rect 13464 2876 15301 2904
rect 13464 2836 13492 2876
rect 15289 2873 15301 2876
rect 15335 2873 15347 2907
rect 15289 2867 15347 2873
rect 16485 2907 16543 2913
rect 16485 2873 16497 2907
rect 16531 2904 16543 2907
rect 16531 2876 19334 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 8312 2808 13492 2836
rect 14093 2839 14151 2845
rect 7837 2799 7895 2805
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 16390 2836 16396 2848
rect 14139 2808 16396 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 17129 2839 17187 2845
rect 17129 2836 17141 2839
rect 16715 2808 17141 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 17129 2805 17141 2808
rect 17175 2805 17187 2839
rect 19306 2836 19334 2876
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19306 2808 19809 2836
rect 17129 2799 17187 2805
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 1104 2746 21436 2768
rect 1104 2694 4338 2746
rect 4390 2694 4402 2746
rect 4454 2694 4466 2746
rect 4518 2694 4530 2746
rect 4582 2694 4594 2746
rect 4646 2694 11116 2746
rect 11168 2694 11180 2746
rect 11232 2694 11244 2746
rect 11296 2694 11308 2746
rect 11360 2694 11372 2746
rect 11424 2694 17893 2746
rect 17945 2694 17957 2746
rect 18009 2694 18021 2746
rect 18073 2694 18085 2746
rect 18137 2694 18149 2746
rect 18201 2694 21436 2746
rect 1104 2672 21436 2694
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 5675 2604 8616 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 4154 2564 4160 2576
rect 2087 2536 4160 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 7009 2567 7067 2573
rect 7009 2533 7021 2567
rect 7055 2564 7067 2567
rect 8478 2564 8484 2576
rect 7055 2536 8484 2564
rect 7055 2533 7067 2536
rect 7009 2527 7067 2533
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 8588 2564 8616 2604
rect 9306 2592 9312 2644
rect 9364 2632 9370 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9364 2604 9505 2632
rect 9364 2592 9370 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 14182 2632 14188 2644
rect 12308 2604 14188 2632
rect 12308 2592 12314 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 16758 2632 16764 2644
rect 14936 2604 16764 2632
rect 11606 2564 11612 2576
rect 8588 2536 11612 2564
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 8996 2468 10425 2496
rect 8996 2456 9002 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10413 2459 10471 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12161 2499 12219 2505
rect 12161 2496 12173 2499
rect 12124 2468 12173 2496
rect 12124 2456 12130 2468
rect 12161 2465 12173 2468
rect 12207 2496 12219 2499
rect 13354 2496 13360 2508
rect 12207 2468 13360 2496
rect 12207 2465 12219 2468
rect 12161 2459 12219 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 1728 2400 2789 2428
rect 1728 2388 1734 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 5350 2388 5356 2440
rect 5408 2428 5414 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5408 2400 5457 2428
rect 5408 2388 5414 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 6512 2400 7757 2428
rect 6512 2388 6518 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 7745 2391 7803 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 14936 2437 14964 2604
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 16899 2635 16957 2641
rect 16899 2601 16911 2635
rect 16945 2632 16957 2635
rect 17678 2632 17684 2644
rect 16945 2604 17684 2632
rect 16945 2601 16957 2604
rect 16899 2595 16957 2601
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 19150 2592 19156 2644
rect 19208 2632 19214 2644
rect 20625 2635 20683 2641
rect 20625 2632 20637 2635
rect 19208 2604 20637 2632
rect 19208 2592 19214 2604
rect 20625 2601 20637 2604
rect 20671 2601 20683 2635
rect 20625 2595 20683 2601
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15841 2567 15899 2573
rect 15841 2564 15853 2567
rect 15620 2536 15853 2564
rect 15620 2524 15626 2536
rect 15841 2533 15853 2536
rect 15887 2533 15899 2567
rect 15841 2527 15899 2533
rect 15105 2499 15163 2505
rect 15105 2465 15117 2499
rect 15151 2496 15163 2499
rect 16942 2496 16948 2508
rect 15151 2468 16948 2496
rect 15151 2465 15163 2468
rect 15105 2459 15163 2465
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 18233 2499 18291 2505
rect 18233 2496 18245 2499
rect 17184 2468 18245 2496
rect 17184 2456 17190 2468
rect 18233 2465 18245 2468
rect 18279 2465 18291 2499
rect 18233 2459 18291 2465
rect 18598 2456 18604 2508
rect 18656 2496 18662 2508
rect 18656 2468 20576 2496
rect 18656 2456 18662 2468
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11848 2400 11897 2428
rect 11848 2388 11854 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16632 2400 16681 2428
rect 16632 2388 16638 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 20548 2437 20576 2468
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19024 2400 19257 2428
rect 19024 2388 19030 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 2464 2332 2605 2360
rect 2464 2320 2470 2332
rect 2593 2329 2605 2332
rect 2639 2329 2651 2363
rect 2593 2323 2651 2329
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 3016 2332 4261 2360
rect 3016 2320 3022 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 6825 2363 6883 2369
rect 6825 2360 6837 2363
rect 5960 2332 6837 2360
rect 5960 2320 5966 2332
rect 6825 2329 6837 2332
rect 6871 2329 6883 2363
rect 6825 2323 6883 2329
rect 7561 2363 7619 2369
rect 7561 2329 7573 2363
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 4338 2292 4344 2304
rect 4299 2264 4344 2292
rect 4338 2252 4344 2264
rect 4396 2252 4402 2304
rect 7576 2292 7604 2323
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 8352 2332 9413 2360
rect 8352 2320 8358 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 12526 2320 12532 2372
rect 12584 2360 12590 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 12584 2332 13277 2360
rect 12584 2320 12590 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 15528 2332 15669 2360
rect 15528 2320 15534 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 17310 2320 17316 2372
rect 17368 2360 17374 2372
rect 18049 2363 18107 2369
rect 18049 2360 18061 2363
rect 17368 2332 18061 2360
rect 17368 2320 17374 2332
rect 18049 2329 18061 2332
rect 18095 2329 18107 2363
rect 18049 2323 18107 2329
rect 13170 2292 13176 2304
rect 7576 2264 13176 2292
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19536 2292 19564 2391
rect 18840 2264 19564 2292
rect 18840 2252 18846 2264
rect 1104 2202 21436 2224
rect 1104 2150 7727 2202
rect 7779 2150 7791 2202
rect 7843 2150 7855 2202
rect 7907 2150 7919 2202
rect 7971 2150 7983 2202
rect 8035 2150 14504 2202
rect 14556 2150 14568 2202
rect 14620 2150 14632 2202
rect 14684 2150 14696 2202
rect 14748 2150 14760 2202
rect 14812 2150 21436 2202
rect 1104 2128 21436 2150
rect 4338 2048 4344 2100
rect 4396 2088 4402 2100
rect 19058 2088 19064 2100
rect 4396 2060 19064 2088
rect 4396 2048 4402 2060
rect 19058 2048 19064 2060
rect 19116 2048 19122 2100
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 13354 2020 13360 2032
rect 7616 1992 13360 2020
rect 7616 1980 7622 1992
rect 13354 1980 13360 1992
rect 13412 1980 13418 2032
rect 16758 1980 16764 2032
rect 16816 2020 16822 2032
rect 19886 2020 19892 2032
rect 16816 1992 19892 2020
rect 16816 1980 16822 1992
rect 19886 1980 19892 1992
rect 19944 1980 19950 2032
<< via1 >>
rect 17868 22448 17920 22500
rect 18328 22448 18380 22500
rect 4338 22278 4390 22330
rect 4402 22278 4454 22330
rect 4466 22278 4518 22330
rect 4530 22278 4582 22330
rect 4594 22278 4646 22330
rect 11116 22278 11168 22330
rect 11180 22278 11232 22330
rect 11244 22278 11296 22330
rect 11308 22278 11360 22330
rect 11372 22278 11424 22330
rect 17893 22278 17945 22330
rect 17957 22278 18009 22330
rect 18021 22278 18073 22330
rect 18085 22278 18137 22330
rect 18149 22278 18201 22330
rect 5356 22108 5408 22160
rect 4068 22040 4120 22092
rect 5724 22040 5776 22092
rect 2780 21972 2832 22024
rect 3516 21972 3568 22024
rect 3608 21904 3660 21956
rect 5908 21972 5960 22024
rect 6276 21972 6328 22024
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6920 22015 6972 22024
rect 6644 21972 6696 21981
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 7564 21972 7616 22024
rect 8300 21972 8352 22024
rect 9956 21972 10008 22024
rect 10600 21972 10652 22024
rect 10876 21972 10928 22024
rect 11152 22040 11204 22092
rect 14832 22176 14884 22228
rect 14740 22040 14792 22092
rect 11704 21972 11756 22024
rect 12440 21972 12492 22024
rect 15384 22040 15436 22092
rect 16856 22040 16908 22092
rect 17408 22040 17460 22092
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 16580 21972 16632 22024
rect 18512 22015 18564 22024
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 21364 22040 21416 22092
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 5540 21836 5592 21888
rect 6000 21836 6052 21888
rect 8944 21836 8996 21888
rect 10508 21836 10560 21888
rect 10876 21879 10928 21888
rect 10876 21845 10885 21879
rect 10885 21845 10919 21879
rect 10919 21845 10928 21879
rect 10876 21836 10928 21845
rect 12164 21836 12216 21888
rect 18972 21904 19024 21956
rect 17040 21836 17092 21888
rect 17224 21836 17276 21888
rect 19340 21836 19392 21888
rect 7727 21734 7779 21786
rect 7791 21734 7843 21786
rect 7855 21734 7907 21786
rect 7919 21734 7971 21786
rect 7983 21734 8035 21786
rect 14504 21734 14556 21786
rect 14568 21734 14620 21786
rect 14632 21734 14684 21786
rect 14696 21734 14748 21786
rect 14760 21734 14812 21786
rect 5356 21632 5408 21684
rect 9404 21632 9456 21684
rect 1860 21607 1912 21616
rect 1860 21573 1869 21607
rect 1869 21573 1903 21607
rect 1903 21573 1912 21607
rect 1860 21564 1912 21573
rect 4896 21564 4948 21616
rect 9312 21564 9364 21616
rect 10232 21632 10284 21684
rect 11520 21632 11572 21684
rect 11428 21564 11480 21616
rect 13728 21632 13780 21684
rect 3148 21496 3200 21548
rect 1768 21360 1820 21412
rect 3056 21292 3108 21344
rect 5448 21496 5500 21548
rect 6184 21496 6236 21548
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 8300 21539 8352 21548
rect 8300 21505 8309 21539
rect 8309 21505 8343 21539
rect 8343 21505 8352 21539
rect 8300 21496 8352 21505
rect 10048 21496 10100 21548
rect 10232 21539 10284 21548
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 5356 21428 5408 21480
rect 6368 21471 6420 21480
rect 6368 21437 6377 21471
rect 6377 21437 6411 21471
rect 6411 21437 6420 21471
rect 6368 21428 6420 21437
rect 7472 21428 7524 21480
rect 8024 21428 8076 21480
rect 7564 21360 7616 21412
rect 8668 21292 8720 21344
rect 9220 21428 9272 21480
rect 11520 21428 11572 21480
rect 12348 21496 12400 21548
rect 13084 21564 13136 21616
rect 13268 21564 13320 21616
rect 13176 21496 13228 21548
rect 13452 21564 13504 21616
rect 13268 21428 13320 21480
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 13820 21496 13872 21548
rect 14832 21632 14884 21684
rect 14464 21564 14516 21616
rect 16028 21564 16080 21616
rect 17040 21632 17092 21684
rect 15016 21539 15068 21548
rect 13636 21428 13688 21480
rect 15016 21505 15025 21539
rect 15025 21505 15059 21539
rect 15059 21505 15068 21539
rect 15016 21496 15068 21505
rect 15844 21496 15896 21548
rect 17500 21496 17552 21548
rect 18236 21496 18288 21548
rect 19064 21496 19116 21548
rect 22468 21496 22520 21548
rect 15292 21428 15344 21480
rect 15476 21428 15528 21480
rect 19432 21428 19484 21480
rect 9128 21360 9180 21412
rect 13176 21360 13228 21412
rect 16580 21360 16632 21412
rect 17408 21360 17460 21412
rect 17592 21360 17644 21412
rect 9956 21292 10008 21344
rect 10324 21292 10376 21344
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 11520 21292 11572 21344
rect 11980 21292 12032 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 12348 21292 12400 21344
rect 12900 21292 12952 21344
rect 15016 21292 15068 21344
rect 15476 21292 15528 21344
rect 17224 21292 17276 21344
rect 17776 21292 17828 21344
rect 18512 21292 18564 21344
rect 4338 21190 4390 21242
rect 4402 21190 4454 21242
rect 4466 21190 4518 21242
rect 4530 21190 4582 21242
rect 4594 21190 4646 21242
rect 11116 21190 11168 21242
rect 11180 21190 11232 21242
rect 11244 21190 11296 21242
rect 11308 21190 11360 21242
rect 11372 21190 11424 21242
rect 17893 21190 17945 21242
rect 17957 21190 18009 21242
rect 18021 21190 18073 21242
rect 18085 21190 18137 21242
rect 18149 21190 18201 21242
rect 572 21088 624 21140
rect 4712 21088 4764 21140
rect 8024 21088 8076 21140
rect 9864 21088 9916 21140
rect 10876 21088 10928 21140
rect 11612 21088 11664 21140
rect 13360 21088 13412 21140
rect 13636 21088 13688 21140
rect 14372 21131 14424 21140
rect 14372 21097 14381 21131
rect 14381 21097 14415 21131
rect 14415 21097 14424 21131
rect 14372 21088 14424 21097
rect 16396 21131 16448 21140
rect 16396 21097 16405 21131
rect 16405 21097 16439 21131
rect 16439 21097 16448 21131
rect 16396 21088 16448 21097
rect 2228 21020 2280 21072
rect 4988 21020 5040 21072
rect 4344 20995 4396 21004
rect 4344 20961 4353 20995
rect 4353 20961 4387 20995
rect 4387 20961 4396 20995
rect 4344 20952 4396 20961
rect 5816 20952 5868 21004
rect 1124 20884 1176 20936
rect 5540 20884 5592 20936
rect 5724 20927 5776 20936
rect 5724 20893 5733 20927
rect 5733 20893 5767 20927
rect 5767 20893 5776 20927
rect 5724 20884 5776 20893
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 7196 21020 7248 21072
rect 8484 20952 8536 21004
rect 2504 20816 2556 20868
rect 4160 20791 4212 20800
rect 4160 20757 4169 20791
rect 4169 20757 4203 20791
rect 4203 20757 4212 20791
rect 4160 20748 4212 20757
rect 4252 20791 4304 20800
rect 4252 20757 4261 20791
rect 4261 20757 4295 20791
rect 4295 20757 4304 20791
rect 5080 20859 5132 20868
rect 5080 20825 5089 20859
rect 5089 20825 5123 20859
rect 5123 20825 5132 20859
rect 5080 20816 5132 20825
rect 6368 20816 6420 20868
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 9220 20927 9272 20936
rect 9220 20893 9229 20927
rect 9229 20893 9263 20927
rect 9263 20893 9272 20927
rect 9220 20884 9272 20893
rect 4252 20748 4304 20757
rect 5540 20748 5592 20800
rect 5632 20748 5684 20800
rect 6276 20791 6328 20800
rect 6276 20757 6285 20791
rect 6285 20757 6319 20791
rect 6319 20757 6328 20791
rect 6276 20748 6328 20757
rect 7656 20748 7708 20800
rect 8116 20816 8168 20868
rect 9128 20748 9180 20800
rect 9588 20952 9640 21004
rect 9772 20952 9824 21004
rect 10416 20952 10468 21004
rect 10784 20952 10836 21004
rect 10140 20884 10192 20936
rect 10324 20927 10376 20936
rect 10324 20893 10333 20927
rect 10333 20893 10367 20927
rect 10367 20893 10376 20927
rect 10324 20884 10376 20893
rect 11060 20952 11112 21004
rect 15844 21020 15896 21072
rect 12532 20952 12584 21004
rect 13820 20952 13872 21004
rect 11980 20884 12032 20936
rect 14004 20884 14056 20936
rect 15108 20884 15160 20936
rect 16120 20952 16172 21004
rect 16948 20952 17000 21004
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 17868 20995 17920 21004
rect 17868 20961 17877 20995
rect 17877 20961 17911 20995
rect 17911 20961 17920 20995
rect 17868 20952 17920 20961
rect 16764 20884 16816 20936
rect 17592 20884 17644 20936
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 19524 20884 19576 20936
rect 21916 20884 21968 20936
rect 10048 20748 10100 20800
rect 13176 20816 13228 20868
rect 13268 20816 13320 20868
rect 13452 20816 13504 20868
rect 14464 20816 14516 20868
rect 15568 20816 15620 20868
rect 17500 20816 17552 20868
rect 11612 20748 11664 20800
rect 12072 20791 12124 20800
rect 12072 20757 12081 20791
rect 12081 20757 12115 20791
rect 12115 20757 12124 20791
rect 12072 20748 12124 20757
rect 12440 20748 12492 20800
rect 13636 20748 13688 20800
rect 13820 20748 13872 20800
rect 14832 20791 14884 20800
rect 14832 20757 14841 20791
rect 14841 20757 14875 20791
rect 14875 20757 14884 20791
rect 14832 20748 14884 20757
rect 16672 20748 16724 20800
rect 17684 20791 17736 20800
rect 17684 20757 17693 20791
rect 17693 20757 17727 20791
rect 17727 20757 17736 20791
rect 17684 20748 17736 20757
rect 19616 20748 19668 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 7727 20646 7779 20698
rect 7791 20646 7843 20698
rect 7855 20646 7907 20698
rect 7919 20646 7971 20698
rect 7983 20646 8035 20698
rect 14504 20646 14556 20698
rect 14568 20646 14620 20698
rect 14632 20646 14684 20698
rect 14696 20646 14748 20698
rect 14760 20646 14812 20698
rect 2320 20587 2372 20596
rect 2320 20553 2329 20587
rect 2329 20553 2363 20587
rect 2363 20553 2372 20587
rect 2320 20544 2372 20553
rect 4160 20544 4212 20596
rect 5356 20544 5408 20596
rect 3056 20476 3108 20528
rect 4252 20476 4304 20528
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 2688 20340 2740 20392
rect 3884 20451 3936 20460
rect 3884 20417 3893 20451
rect 3893 20417 3927 20451
rect 3927 20417 3936 20451
rect 3884 20408 3936 20417
rect 4804 20408 4856 20460
rect 5908 20544 5960 20596
rect 6920 20544 6972 20596
rect 8116 20544 8168 20596
rect 8668 20587 8720 20596
rect 8668 20553 8677 20587
rect 8677 20553 8711 20587
rect 8711 20553 8720 20587
rect 8668 20544 8720 20553
rect 9772 20544 9824 20596
rect 10232 20544 10284 20596
rect 10416 20544 10468 20596
rect 10876 20544 10928 20596
rect 11520 20544 11572 20596
rect 6276 20476 6328 20528
rect 7288 20476 7340 20528
rect 7380 20476 7432 20528
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6092 20408 6144 20460
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 6644 20408 6696 20417
rect 7656 20451 7708 20460
rect 2872 20272 2924 20324
rect 5356 20340 5408 20392
rect 6276 20340 6328 20392
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8392 20476 8444 20528
rect 8208 20451 8260 20460
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 8668 20451 8720 20460
rect 8668 20417 8677 20451
rect 8677 20417 8711 20451
rect 8711 20417 8720 20451
rect 8668 20408 8720 20417
rect 8760 20408 8812 20460
rect 9680 20476 9732 20528
rect 9864 20451 9916 20460
rect 7012 20340 7064 20392
rect 7748 20340 7800 20392
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 11612 20451 11664 20460
rect 11612 20417 11621 20451
rect 11621 20417 11655 20451
rect 11655 20417 11664 20451
rect 11612 20408 11664 20417
rect 10692 20383 10744 20392
rect 10692 20349 10701 20383
rect 10701 20349 10735 20383
rect 10735 20349 10744 20383
rect 10692 20340 10744 20349
rect 14188 20476 14240 20528
rect 14832 20544 14884 20596
rect 15108 20544 15160 20596
rect 16580 20544 16632 20596
rect 17684 20587 17736 20596
rect 17684 20553 17693 20587
rect 17693 20553 17727 20587
rect 17727 20553 17736 20587
rect 17684 20544 17736 20553
rect 19248 20544 19300 20596
rect 16212 20476 16264 20528
rect 11980 20408 12032 20460
rect 12440 20408 12492 20460
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 13268 20451 13320 20460
rect 12992 20408 13044 20417
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 14372 20408 14424 20460
rect 14832 20451 14884 20460
rect 14832 20417 14841 20451
rect 14841 20417 14875 20451
rect 14875 20417 14884 20451
rect 15108 20451 15160 20460
rect 14832 20408 14884 20417
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 15292 20408 15344 20460
rect 5448 20272 5500 20324
rect 6184 20272 6236 20324
rect 8300 20272 8352 20324
rect 9588 20272 9640 20324
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 3976 20204 4028 20256
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 6828 20204 6880 20256
rect 7472 20204 7524 20256
rect 7656 20204 7708 20256
rect 8576 20204 8628 20256
rect 9956 20204 10008 20256
rect 10232 20272 10284 20324
rect 10968 20204 11020 20256
rect 15660 20340 15712 20392
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 16396 20408 16448 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 17316 20476 17368 20528
rect 18512 20476 18564 20528
rect 20260 20476 20312 20528
rect 16304 20340 16356 20392
rect 18788 20451 18840 20460
rect 18788 20417 18797 20451
rect 18797 20417 18831 20451
rect 18831 20417 18840 20451
rect 18788 20408 18840 20417
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 17592 20340 17644 20392
rect 13176 20315 13228 20324
rect 13176 20281 13185 20315
rect 13185 20281 13219 20315
rect 13219 20281 13228 20315
rect 13176 20272 13228 20281
rect 13360 20272 13412 20324
rect 15016 20247 15068 20256
rect 15016 20213 15025 20247
rect 15025 20213 15059 20247
rect 15059 20213 15068 20247
rect 15016 20204 15068 20213
rect 15752 20204 15804 20256
rect 16580 20204 16632 20256
rect 18972 20247 19024 20256
rect 18972 20213 18981 20247
rect 18981 20213 19015 20247
rect 19015 20213 19024 20247
rect 18972 20204 19024 20213
rect 20076 20204 20128 20256
rect 4338 20102 4390 20154
rect 4402 20102 4454 20154
rect 4466 20102 4518 20154
rect 4530 20102 4582 20154
rect 4594 20102 4646 20154
rect 11116 20102 11168 20154
rect 11180 20102 11232 20154
rect 11244 20102 11296 20154
rect 11308 20102 11360 20154
rect 11372 20102 11424 20154
rect 17893 20102 17945 20154
rect 17957 20102 18009 20154
rect 18021 20102 18073 20154
rect 18085 20102 18137 20154
rect 18149 20102 18201 20154
rect 4712 20000 4764 20052
rect 6460 20043 6512 20052
rect 1676 19932 1728 19984
rect 5908 19932 5960 19984
rect 6460 20009 6469 20043
rect 6469 20009 6503 20043
rect 6503 20009 6512 20043
rect 6460 20000 6512 20009
rect 8668 20000 8720 20052
rect 8852 20000 8904 20052
rect 13728 20000 13780 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 16028 20000 16080 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 17132 20043 17184 20052
rect 17132 20009 17141 20043
rect 17141 20009 17175 20043
rect 17175 20009 17184 20043
rect 17132 20000 17184 20009
rect 18420 20000 18472 20052
rect 8208 19932 8260 19984
rect 11520 19932 11572 19984
rect 4344 19907 4396 19916
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 4344 19873 4353 19907
rect 4353 19873 4387 19907
rect 4387 19873 4396 19907
rect 4344 19864 4396 19873
rect 4528 19864 4580 19916
rect 7012 19864 7064 19916
rect 7196 19864 7248 19916
rect 7656 19864 7708 19916
rect 8116 19864 8168 19916
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 10048 19864 10100 19916
rect 10784 19864 10836 19916
rect 11796 19932 11848 19984
rect 18328 19932 18380 19984
rect 4712 19796 4764 19848
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 5448 19796 5500 19805
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 7748 19839 7800 19848
rect 2872 19771 2924 19780
rect 2872 19737 2881 19771
rect 2881 19737 2915 19771
rect 2915 19737 2924 19771
rect 2872 19728 2924 19737
rect 3056 19771 3108 19780
rect 3056 19737 3065 19771
rect 3065 19737 3099 19771
rect 3099 19737 3108 19771
rect 3056 19728 3108 19737
rect 3148 19660 3200 19712
rect 4068 19660 4120 19712
rect 4252 19703 4304 19712
rect 4252 19669 4261 19703
rect 4261 19669 4295 19703
rect 4295 19669 4304 19703
rect 4252 19660 4304 19669
rect 5172 19660 5224 19712
rect 5632 19660 5684 19712
rect 5816 19703 5868 19712
rect 5816 19669 5825 19703
rect 5825 19669 5859 19703
rect 5859 19669 5868 19703
rect 5816 19660 5868 19669
rect 6736 19728 6788 19780
rect 7748 19805 7757 19839
rect 7757 19805 7791 19839
rect 7791 19805 7800 19839
rect 7748 19796 7800 19805
rect 7840 19796 7892 19848
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 8668 19796 8720 19848
rect 9312 19796 9364 19848
rect 9588 19796 9640 19848
rect 12716 19796 12768 19848
rect 8116 19728 8168 19780
rect 8484 19728 8536 19780
rect 9036 19728 9088 19780
rect 10876 19728 10928 19780
rect 18236 19864 18288 19916
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 15476 19796 15528 19848
rect 15844 19796 15896 19848
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 17224 19796 17276 19848
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 14096 19728 14148 19780
rect 15936 19728 15988 19780
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 18604 19728 18656 19780
rect 19800 19771 19852 19780
rect 19800 19737 19809 19771
rect 19809 19737 19843 19771
rect 19843 19737 19852 19771
rect 19800 19728 19852 19737
rect 9680 19660 9732 19712
rect 9864 19703 9916 19712
rect 9864 19669 9873 19703
rect 9873 19669 9907 19703
rect 9907 19669 9916 19703
rect 9864 19660 9916 19669
rect 11980 19660 12032 19712
rect 12348 19703 12400 19712
rect 12348 19669 12357 19703
rect 12357 19669 12391 19703
rect 12391 19669 12400 19703
rect 12348 19660 12400 19669
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 12716 19660 12768 19669
rect 15660 19660 15712 19712
rect 16488 19660 16540 19712
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 7727 19558 7779 19610
rect 7791 19558 7843 19610
rect 7855 19558 7907 19610
rect 7919 19558 7971 19610
rect 7983 19558 8035 19610
rect 14504 19558 14556 19610
rect 14568 19558 14620 19610
rect 14632 19558 14684 19610
rect 14696 19558 14748 19610
rect 14760 19558 14812 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 3148 19456 3200 19508
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 5724 19456 5776 19508
rect 3884 19388 3936 19440
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 1216 19252 1268 19304
rect 1676 19320 1728 19372
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 4528 19363 4580 19372
rect 4528 19329 4537 19363
rect 4537 19329 4571 19363
rect 4571 19329 4580 19363
rect 4528 19320 4580 19329
rect 4988 19363 5040 19372
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 2872 19252 2924 19304
rect 3056 19252 3108 19304
rect 3792 19252 3844 19304
rect 4160 19252 4212 19304
rect 5908 19388 5960 19440
rect 6276 19388 6328 19440
rect 8668 19456 8720 19508
rect 9864 19456 9916 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 13728 19456 13780 19508
rect 7012 19388 7064 19440
rect 8484 19388 8536 19440
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 7288 19320 7340 19372
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 8760 19320 8812 19372
rect 9128 19320 9180 19372
rect 9312 19320 9364 19372
rect 9772 19320 9824 19372
rect 9956 19363 10008 19372
rect 9956 19329 9965 19363
rect 9965 19329 9999 19363
rect 9999 19329 10008 19363
rect 9956 19320 10008 19329
rect 10140 19363 10192 19372
rect 10140 19329 10149 19363
rect 10149 19329 10183 19363
rect 10183 19329 10192 19363
rect 10140 19320 10192 19329
rect 10232 19363 10284 19372
rect 10232 19329 10241 19363
rect 10241 19329 10275 19363
rect 10275 19329 10284 19363
rect 11704 19388 11756 19440
rect 10232 19320 10284 19329
rect 10600 19320 10652 19372
rect 11980 19363 12032 19372
rect 11980 19329 11989 19363
rect 11989 19329 12023 19363
rect 12023 19329 12032 19363
rect 11980 19320 12032 19329
rect 12072 19320 12124 19372
rect 12716 19388 12768 19440
rect 12808 19388 12860 19440
rect 13360 19388 13412 19440
rect 14004 19431 14056 19440
rect 14004 19397 14013 19431
rect 14013 19397 14047 19431
rect 14047 19397 14056 19431
rect 14004 19388 14056 19397
rect 10968 19252 11020 19304
rect 11520 19252 11572 19304
rect 13176 19320 13228 19372
rect 15752 19456 15804 19508
rect 16304 19456 16356 19508
rect 13820 19252 13872 19304
rect 14188 19320 14240 19372
rect 15476 19320 15528 19372
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 16028 19363 16080 19372
rect 15844 19320 15896 19329
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 17500 19388 17552 19440
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 19340 19388 19392 19440
rect 18512 19320 18564 19372
rect 19248 19320 19300 19372
rect 3884 19184 3936 19236
rect 5540 19184 5592 19236
rect 6184 19184 6236 19236
rect 12440 19184 12492 19236
rect 12992 19184 13044 19236
rect 15844 19184 15896 19236
rect 18328 19252 18380 19304
rect 18972 19252 19024 19304
rect 19156 19252 19208 19304
rect 20812 19184 20864 19236
rect 4068 19116 4120 19168
rect 6092 19116 6144 19168
rect 7104 19116 7156 19168
rect 10232 19116 10284 19168
rect 12256 19116 12308 19168
rect 14188 19116 14240 19168
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15660 19116 15712 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 18236 19116 18288 19168
rect 4338 19014 4390 19066
rect 4402 19014 4454 19066
rect 4466 19014 4518 19066
rect 4530 19014 4582 19066
rect 4594 19014 4646 19066
rect 11116 19014 11168 19066
rect 11180 19014 11232 19066
rect 11244 19014 11296 19066
rect 11308 19014 11360 19066
rect 11372 19014 11424 19066
rect 17893 19014 17945 19066
rect 17957 19014 18009 19066
rect 18021 19014 18073 19066
rect 18085 19014 18137 19066
rect 18149 19014 18201 19066
rect 2228 18912 2280 18964
rect 2964 18912 3016 18964
rect 4160 18912 4212 18964
rect 5172 18912 5224 18964
rect 6644 18912 6696 18964
rect 9036 18912 9088 18964
rect 11980 18912 12032 18964
rect 14188 18955 14240 18964
rect 14188 18921 14197 18955
rect 14197 18921 14231 18955
rect 14231 18921 14240 18955
rect 14188 18912 14240 18921
rect 14924 18912 14976 18964
rect 16764 18955 16816 18964
rect 2228 18819 2280 18828
rect 2228 18785 2237 18819
rect 2237 18785 2271 18819
rect 2271 18785 2280 18819
rect 2228 18776 2280 18785
rect 5816 18776 5868 18828
rect 6368 18776 6420 18828
rect 6736 18844 6788 18896
rect 10324 18844 10376 18896
rect 7288 18776 7340 18828
rect 11520 18844 11572 18896
rect 13360 18844 13412 18896
rect 2136 18708 2188 18760
rect 2596 18708 2648 18760
rect 3792 18751 3844 18760
rect 3792 18717 3801 18751
rect 3801 18717 3835 18751
rect 3835 18717 3844 18751
rect 3792 18708 3844 18717
rect 3884 18708 3936 18760
rect 5448 18640 5500 18692
rect 5908 18708 5960 18760
rect 6736 18708 6788 18760
rect 5816 18640 5868 18692
rect 7196 18708 7248 18760
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 9036 18708 9088 18717
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 10784 18776 10836 18828
rect 10876 18708 10928 18760
rect 12072 18776 12124 18828
rect 13176 18819 13228 18828
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 10140 18640 10192 18692
rect 12348 18708 12400 18760
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 12072 18640 12124 18692
rect 14004 18708 14056 18760
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 16764 18921 16773 18955
rect 16773 18921 16807 18955
rect 16807 18921 16816 18955
rect 16764 18912 16816 18921
rect 16948 18912 17000 18964
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 16488 18751 16540 18760
rect 15844 18708 15896 18717
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 16672 18844 16724 18896
rect 17776 18912 17828 18964
rect 19800 18912 19852 18964
rect 17592 18776 17644 18828
rect 20628 18776 20680 18828
rect 16764 18708 16816 18760
rect 18236 18708 18288 18760
rect 18420 18708 18472 18760
rect 18788 18708 18840 18760
rect 15108 18640 15160 18692
rect 19800 18640 19852 18692
rect 3424 18572 3476 18624
rect 5632 18572 5684 18624
rect 5724 18572 5776 18624
rect 6184 18572 6236 18624
rect 6920 18572 6972 18624
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 12256 18572 12308 18624
rect 12900 18572 12952 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 14280 18572 14332 18624
rect 14924 18572 14976 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 19340 18572 19392 18624
rect 7727 18470 7779 18522
rect 7791 18470 7843 18522
rect 7855 18470 7907 18522
rect 7919 18470 7971 18522
rect 7983 18470 8035 18522
rect 14504 18470 14556 18522
rect 14568 18470 14620 18522
rect 14632 18470 14684 18522
rect 14696 18470 14748 18522
rect 14760 18470 14812 18522
rect 1676 18411 1728 18420
rect 1676 18377 1685 18411
rect 1685 18377 1719 18411
rect 1719 18377 1728 18411
rect 1676 18368 1728 18377
rect 2596 18411 2648 18420
rect 2596 18377 2605 18411
rect 2605 18377 2639 18411
rect 2639 18377 2648 18411
rect 2596 18368 2648 18377
rect 3424 18411 3476 18420
rect 3424 18377 3433 18411
rect 3433 18377 3467 18411
rect 3467 18377 3476 18411
rect 3424 18368 3476 18377
rect 2412 18343 2464 18352
rect 2412 18309 2421 18343
rect 2421 18309 2455 18343
rect 2455 18309 2464 18343
rect 2412 18300 2464 18309
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 5724 18368 5776 18420
rect 6552 18368 6604 18420
rect 7012 18411 7064 18420
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 10324 18368 10376 18420
rect 12992 18368 13044 18420
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 15660 18368 15712 18420
rect 16120 18368 16172 18420
rect 17684 18368 17736 18420
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 20260 18368 20312 18420
rect 7196 18300 7248 18352
rect 7288 18300 7340 18352
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 3976 18232 4028 18284
rect 5080 18232 5132 18284
rect 5356 18232 5408 18284
rect 5632 18275 5684 18284
rect 3332 18164 3384 18216
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 6368 18275 6420 18284
rect 6368 18241 6377 18275
rect 6377 18241 6411 18275
rect 6411 18241 6420 18275
rect 6368 18232 6420 18241
rect 6644 18275 6696 18284
rect 6644 18241 6653 18275
rect 6653 18241 6687 18275
rect 6687 18241 6696 18275
rect 6644 18232 6696 18241
rect 6552 18164 6604 18216
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 8576 18232 8628 18284
rect 9128 18232 9180 18284
rect 9220 18232 9272 18284
rect 10324 18232 10376 18284
rect 10692 18232 10744 18284
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11980 18232 12032 18284
rect 12532 18232 12584 18284
rect 8760 18164 8812 18216
rect 9772 18207 9824 18216
rect 9772 18173 9781 18207
rect 9781 18173 9815 18207
rect 9815 18173 9824 18207
rect 9772 18164 9824 18173
rect 10048 18164 10100 18216
rect 5540 18096 5592 18148
rect 5632 18096 5684 18148
rect 6736 18096 6788 18148
rect 12072 18096 12124 18148
rect 12624 18096 12676 18148
rect 12900 18232 12952 18284
rect 13176 18232 13228 18284
rect 13820 18232 13872 18284
rect 15108 18232 15160 18284
rect 16028 18232 16080 18284
rect 16212 18300 16264 18352
rect 16580 18232 16632 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 17776 18232 17828 18284
rect 18788 18232 18840 18284
rect 19064 18275 19116 18284
rect 19064 18241 19073 18275
rect 19073 18241 19107 18275
rect 19107 18241 19116 18275
rect 19064 18232 19116 18241
rect 19984 18275 20036 18284
rect 19984 18241 19990 18275
rect 19990 18241 20024 18275
rect 20024 18241 20036 18275
rect 19984 18232 20036 18241
rect 15476 18164 15528 18216
rect 15752 18164 15804 18216
rect 16764 18164 16816 18216
rect 14188 18096 14240 18148
rect 4252 18028 4304 18080
rect 7012 18028 7064 18080
rect 13084 18028 13136 18080
rect 13268 18028 13320 18080
rect 18696 18096 18748 18148
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 15660 18028 15712 18080
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 16028 18028 16080 18080
rect 16396 18028 16448 18080
rect 17040 18028 17092 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 18972 18028 19024 18080
rect 20260 18028 20312 18080
rect 4338 17926 4390 17978
rect 4402 17926 4454 17978
rect 4466 17926 4518 17978
rect 4530 17926 4582 17978
rect 4594 17926 4646 17978
rect 11116 17926 11168 17978
rect 11180 17926 11232 17978
rect 11244 17926 11296 17978
rect 11308 17926 11360 17978
rect 11372 17926 11424 17978
rect 17893 17926 17945 17978
rect 17957 17926 18009 17978
rect 18021 17926 18073 17978
rect 18085 17926 18137 17978
rect 18149 17926 18201 17978
rect 5724 17824 5776 17876
rect 6552 17824 6604 17876
rect 9220 17824 9272 17876
rect 9496 17824 9548 17876
rect 10692 17824 10744 17876
rect 12072 17867 12124 17876
rect 12072 17833 12081 17867
rect 12081 17833 12115 17867
rect 12115 17833 12124 17867
rect 12072 17824 12124 17833
rect 12624 17824 12676 17876
rect 13728 17824 13780 17876
rect 14280 17824 14332 17876
rect 14832 17824 14884 17876
rect 15568 17824 15620 17876
rect 16028 17824 16080 17876
rect 16304 17824 16356 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 19340 17824 19392 17876
rect 2412 17688 2464 17740
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3976 17688 4028 17740
rect 4160 17688 4212 17740
rect 5264 17756 5316 17808
rect 7840 17756 7892 17808
rect 9036 17756 9088 17808
rect 9956 17799 10008 17808
rect 3332 17620 3384 17672
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5816 17620 5868 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 8668 17688 8720 17740
rect 9128 17688 9180 17740
rect 9956 17765 9965 17799
rect 9965 17765 9999 17799
rect 9999 17765 10008 17799
rect 9956 17756 10008 17765
rect 18420 17756 18472 17808
rect 19524 17756 19576 17808
rect 20444 17756 20496 17808
rect 1860 17595 1912 17604
rect 1860 17561 1869 17595
rect 1869 17561 1903 17595
rect 1903 17561 1912 17595
rect 1860 17552 1912 17561
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 3884 17484 3936 17536
rect 4160 17527 4212 17536
rect 4160 17493 4169 17527
rect 4169 17493 4203 17527
rect 4203 17493 4212 17527
rect 4160 17484 4212 17493
rect 5080 17527 5132 17536
rect 5080 17493 5089 17527
rect 5089 17493 5123 17527
rect 5123 17493 5132 17527
rect 5080 17484 5132 17493
rect 6644 17620 6696 17672
rect 6736 17620 6788 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7564 17620 7616 17672
rect 8484 17620 8536 17672
rect 8760 17620 8812 17672
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 9496 17663 9548 17672
rect 6828 17552 6880 17604
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 10140 17620 10192 17672
rect 10324 17620 10376 17672
rect 10692 17620 10744 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 8484 17484 8536 17536
rect 10232 17552 10284 17604
rect 10600 17552 10652 17604
rect 12440 17688 12492 17740
rect 12716 17688 12768 17740
rect 14004 17688 14056 17740
rect 12532 17620 12584 17672
rect 13636 17620 13688 17672
rect 13820 17620 13872 17672
rect 14924 17688 14976 17740
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 16580 17688 16632 17740
rect 17132 17688 17184 17740
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15384 17620 15436 17672
rect 9312 17484 9364 17536
rect 12440 17484 12492 17536
rect 15568 17552 15620 17604
rect 16028 17620 16080 17672
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16488 17552 16540 17604
rect 16948 17620 17000 17672
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18696 17663 18748 17672
rect 18420 17620 18472 17629
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 19984 17620 20036 17672
rect 20536 17663 20588 17672
rect 17776 17484 17828 17536
rect 18788 17552 18840 17604
rect 19340 17552 19392 17604
rect 20536 17629 20545 17663
rect 20545 17629 20579 17663
rect 20579 17629 20588 17663
rect 20536 17620 20588 17629
rect 20628 17620 20680 17672
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 7727 17382 7779 17434
rect 7791 17382 7843 17434
rect 7855 17382 7907 17434
rect 7919 17382 7971 17434
rect 7983 17382 8035 17434
rect 14504 17382 14556 17434
rect 14568 17382 14620 17434
rect 14632 17382 14684 17434
rect 14696 17382 14748 17434
rect 14760 17382 14812 17434
rect 1584 17280 1636 17332
rect 2504 17323 2556 17332
rect 2504 17289 2513 17323
rect 2513 17289 2547 17323
rect 2547 17289 2556 17323
rect 2504 17280 2556 17289
rect 4160 17280 4212 17332
rect 5080 17280 5132 17332
rect 6552 17323 6604 17332
rect 2044 17144 2096 17196
rect 5540 17212 5592 17264
rect 3700 17144 3752 17196
rect 4252 17144 4304 17196
rect 6552 17289 6561 17323
rect 6561 17289 6595 17323
rect 6595 17289 6604 17323
rect 6552 17280 6604 17289
rect 7012 17280 7064 17332
rect 6184 17212 6236 17264
rect 4068 17008 4120 17060
rect 5172 17076 5224 17128
rect 6828 17144 6880 17196
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 5816 17076 5868 17128
rect 8300 17212 8352 17264
rect 8760 17212 8812 17264
rect 9772 17280 9824 17332
rect 11336 17280 11388 17332
rect 13268 17280 13320 17332
rect 13452 17280 13504 17332
rect 14004 17280 14056 17332
rect 14280 17280 14332 17332
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 14832 17280 14884 17332
rect 20076 17280 20128 17332
rect 20260 17323 20312 17332
rect 20260 17289 20269 17323
rect 20269 17289 20303 17323
rect 20303 17289 20312 17323
rect 20260 17280 20312 17289
rect 20628 17323 20680 17332
rect 20628 17289 20637 17323
rect 20637 17289 20671 17323
rect 20671 17289 20680 17323
rect 20628 17280 20680 17289
rect 8668 17187 8720 17196
rect 7380 17076 7432 17128
rect 7472 17076 7524 17128
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 8852 17076 8904 17128
rect 11980 17212 12032 17264
rect 10600 17144 10652 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10876 17144 10928 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 19432 17212 19484 17264
rect 12072 17076 12124 17128
rect 14188 17144 14240 17196
rect 15292 17144 15344 17196
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15568 17187 15620 17196
rect 15384 17144 15436 17153
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 15936 17144 15988 17196
rect 16580 17144 16632 17196
rect 17500 17144 17552 17196
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 18512 17144 18564 17196
rect 18880 17144 18932 17196
rect 19708 17144 19760 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 20536 17144 20588 17196
rect 13176 17076 13228 17128
rect 16672 17076 16724 17128
rect 17132 17076 17184 17128
rect 14004 17008 14056 17060
rect 18144 17076 18196 17128
rect 18696 17076 18748 17128
rect 18788 17051 18840 17060
rect 18788 17017 18797 17051
rect 18797 17017 18831 17051
rect 18831 17017 18840 17051
rect 18788 17008 18840 17017
rect 6368 16940 6420 16992
rect 7104 16940 7156 16992
rect 8668 16940 8720 16992
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 9772 16940 9824 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 12348 16983 12400 16992
rect 12348 16949 12357 16983
rect 12357 16949 12391 16983
rect 12391 16949 12400 16983
rect 12348 16940 12400 16949
rect 12440 16940 12492 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 18880 16940 18932 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 20076 16940 20128 16992
rect 4338 16838 4390 16890
rect 4402 16838 4454 16890
rect 4466 16838 4518 16890
rect 4530 16838 4582 16890
rect 4594 16838 4646 16890
rect 11116 16838 11168 16890
rect 11180 16838 11232 16890
rect 11244 16838 11296 16890
rect 11308 16838 11360 16890
rect 11372 16838 11424 16890
rect 17893 16838 17945 16890
rect 17957 16838 18009 16890
rect 18021 16838 18073 16890
rect 18085 16838 18137 16890
rect 18149 16838 18201 16890
rect 4988 16736 5040 16788
rect 5172 16736 5224 16788
rect 7196 16736 7248 16788
rect 7380 16736 7432 16788
rect 9220 16736 9272 16788
rect 14188 16736 14240 16788
rect 14372 16779 14424 16788
rect 14372 16745 14381 16779
rect 14381 16745 14415 16779
rect 14415 16745 14424 16779
rect 14372 16736 14424 16745
rect 15292 16736 15344 16788
rect 16120 16736 16172 16788
rect 16764 16736 16816 16788
rect 17224 16736 17276 16788
rect 19616 16736 19668 16788
rect 1308 16532 1360 16584
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2780 16532 2832 16584
rect 3240 16532 3292 16584
rect 6828 16668 6880 16720
rect 4252 16532 4304 16584
rect 4712 16532 4764 16584
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 8852 16668 8904 16720
rect 13728 16668 13780 16720
rect 14004 16668 14056 16720
rect 18052 16668 18104 16720
rect 5356 16600 5408 16609
rect 3884 16464 3936 16516
rect 7012 16532 7064 16584
rect 7288 16532 7340 16584
rect 7472 16532 7524 16584
rect 9312 16600 9364 16652
rect 10232 16600 10284 16652
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 12072 16600 12124 16652
rect 12716 16600 12768 16652
rect 14372 16600 14424 16652
rect 11704 16532 11756 16584
rect 13636 16532 13688 16584
rect 14280 16575 14332 16584
rect 7380 16464 7432 16516
rect 2688 16439 2740 16448
rect 2688 16405 2697 16439
rect 2697 16405 2731 16439
rect 2731 16405 2740 16439
rect 2688 16396 2740 16405
rect 4068 16396 4120 16448
rect 4896 16396 4948 16448
rect 5724 16396 5776 16448
rect 7196 16396 7248 16448
rect 8116 16464 8168 16516
rect 9680 16464 9732 16516
rect 7656 16396 7708 16448
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 10968 16396 11020 16448
rect 11980 16396 12032 16448
rect 13912 16464 13964 16516
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16488 16600 16540 16652
rect 19708 16668 19760 16720
rect 20352 16600 20404 16652
rect 15384 16532 15436 16584
rect 14924 16464 14976 16516
rect 15936 16532 15988 16584
rect 16396 16532 16448 16584
rect 16764 16532 16816 16584
rect 17040 16532 17092 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18052 16532 18104 16584
rect 18512 16532 18564 16584
rect 18788 16532 18840 16584
rect 19340 16532 19392 16584
rect 15476 16396 15528 16448
rect 16580 16396 16632 16448
rect 17132 16396 17184 16448
rect 17684 16439 17736 16448
rect 17684 16405 17693 16439
rect 17693 16405 17727 16439
rect 17727 16405 17736 16439
rect 17684 16396 17736 16405
rect 18880 16396 18932 16448
rect 7727 16294 7779 16346
rect 7791 16294 7843 16346
rect 7855 16294 7907 16346
rect 7919 16294 7971 16346
rect 7983 16294 8035 16346
rect 14504 16294 14556 16346
rect 14568 16294 14620 16346
rect 14632 16294 14684 16346
rect 14696 16294 14748 16346
rect 14760 16294 14812 16346
rect 1492 16192 1544 16244
rect 3792 16192 3844 16244
rect 4988 16192 5040 16244
rect 6276 16192 6328 16244
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 10232 16192 10284 16244
rect 13268 16192 13320 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 15476 16192 15528 16244
rect 17684 16235 17736 16244
rect 6368 16124 6420 16176
rect 8392 16124 8444 16176
rect 10048 16124 10100 16176
rect 12992 16124 13044 16176
rect 14280 16124 14332 16176
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 3792 16056 3844 16108
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 2228 16031 2280 16040
rect 2228 15997 2237 16031
rect 2237 15997 2271 16031
rect 2271 15997 2280 16031
rect 2228 15988 2280 15997
rect 2872 15988 2924 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 7656 16056 7708 16108
rect 10416 16056 10468 16108
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 13820 16056 13872 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 15016 16124 15068 16176
rect 5816 15988 5868 16040
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 4160 15920 4212 15972
rect 4896 15963 4948 15972
rect 4896 15929 4905 15963
rect 4905 15929 4939 15963
rect 4939 15929 4948 15963
rect 4896 15920 4948 15929
rect 6828 15988 6880 16040
rect 10784 15988 10836 16040
rect 11520 15988 11572 16040
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 12348 16031 12400 16040
rect 12348 15997 12357 16031
rect 12357 15997 12391 16031
rect 12391 15997 12400 16031
rect 12348 15988 12400 15997
rect 8208 15920 8260 15972
rect 6736 15895 6788 15904
rect 6736 15861 6745 15895
rect 6745 15861 6779 15895
rect 6779 15861 6788 15895
rect 6736 15852 6788 15861
rect 9864 15852 9916 15904
rect 10048 15852 10100 15904
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 13636 15920 13688 15972
rect 13820 15852 13872 15904
rect 14096 15852 14148 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 15568 15920 15620 15972
rect 15752 16056 15804 16108
rect 16580 16056 16632 16108
rect 17684 16201 17693 16235
rect 17693 16201 17727 16235
rect 17727 16201 17736 16235
rect 17684 16192 17736 16201
rect 17132 16124 17184 16176
rect 18604 16056 18656 16108
rect 19248 16056 19300 16108
rect 20536 16056 20588 16108
rect 17040 15988 17092 16040
rect 17592 15988 17644 16040
rect 17684 15920 17736 15972
rect 18788 15988 18840 16040
rect 20260 16031 20312 16040
rect 19248 15920 19300 15972
rect 20260 15997 20269 16031
rect 20269 15997 20303 16031
rect 20303 15997 20312 16031
rect 20260 15988 20312 15997
rect 20720 15920 20772 15972
rect 15660 15852 15712 15904
rect 16212 15852 16264 15904
rect 16672 15852 16724 15904
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 4338 15750 4390 15802
rect 4402 15750 4454 15802
rect 4466 15750 4518 15802
rect 4530 15750 4582 15802
rect 4594 15750 4646 15802
rect 11116 15750 11168 15802
rect 11180 15750 11232 15802
rect 11244 15750 11296 15802
rect 11308 15750 11360 15802
rect 11372 15750 11424 15802
rect 17893 15750 17945 15802
rect 17957 15750 18009 15802
rect 18021 15750 18073 15802
rect 18085 15750 18137 15802
rect 18149 15750 18201 15802
rect 2044 15648 2096 15700
rect 3792 15648 3844 15700
rect 8484 15648 8536 15700
rect 9036 15648 9088 15700
rect 9680 15648 9732 15700
rect 1768 15580 1820 15632
rect 3976 15580 4028 15632
rect 2596 15512 2648 15564
rect 5264 15580 5316 15632
rect 4988 15512 5040 15564
rect 6552 15580 6604 15632
rect 10048 15580 10100 15632
rect 7104 15512 7156 15564
rect 7564 15512 7616 15564
rect 9404 15512 9456 15564
rect 9588 15512 9640 15564
rect 10600 15512 10652 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2688 15444 2740 15496
rect 2780 15444 2832 15496
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 2504 15376 2556 15428
rect 5724 15444 5776 15496
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 9956 15444 10008 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11980 15648 12032 15700
rect 14556 15648 14608 15700
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 17592 15691 17644 15700
rect 17592 15657 17601 15691
rect 17601 15657 17635 15691
rect 17635 15657 17644 15691
rect 17592 15648 17644 15657
rect 18696 15648 18748 15700
rect 3240 15308 3292 15360
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 5724 15351 5776 15360
rect 4620 15308 4672 15317
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 6552 15308 6604 15360
rect 8300 15308 8352 15360
rect 10784 15376 10836 15428
rect 11796 15580 11848 15632
rect 12348 15580 12400 15632
rect 12900 15512 12952 15564
rect 14832 15512 14884 15564
rect 11980 15444 12032 15496
rect 12808 15444 12860 15496
rect 13636 15444 13688 15496
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 16672 15512 16724 15564
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16120 15444 16172 15496
rect 11336 15376 11388 15428
rect 12900 15419 12952 15428
rect 12900 15385 12909 15419
rect 12909 15385 12943 15419
rect 12943 15385 12952 15419
rect 12900 15376 12952 15385
rect 14924 15376 14976 15428
rect 17592 15419 17644 15428
rect 17592 15385 17601 15419
rect 17601 15385 17635 15419
rect 17635 15385 17644 15419
rect 17592 15376 17644 15385
rect 9036 15308 9088 15360
rect 11888 15308 11940 15360
rect 12256 15308 12308 15360
rect 12532 15308 12584 15360
rect 14280 15308 14332 15360
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 18328 15444 18380 15496
rect 18880 15444 18932 15496
rect 19156 15444 19208 15496
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 18236 15308 18288 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 7727 15206 7779 15258
rect 7791 15206 7843 15258
rect 7855 15206 7907 15258
rect 7919 15206 7971 15258
rect 7983 15206 8035 15258
rect 14504 15206 14556 15258
rect 14568 15206 14620 15258
rect 14632 15206 14684 15258
rect 14696 15206 14748 15258
rect 14760 15206 14812 15258
rect 2964 15104 3016 15156
rect 4804 15104 4856 15156
rect 5724 15104 5776 15156
rect 7656 15104 7708 15156
rect 9956 15104 10008 15156
rect 10692 15104 10744 15156
rect 12256 15104 12308 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 15568 15104 15620 15156
rect 16028 15104 16080 15156
rect 17500 15104 17552 15156
rect 20076 15104 20128 15156
rect 20444 15104 20496 15156
rect 3240 15079 3292 15088
rect 2596 14968 2648 15020
rect 3240 15045 3249 15079
rect 3249 15045 3283 15079
rect 3283 15045 3292 15079
rect 3240 15036 3292 15045
rect 4896 15036 4948 15088
rect 4988 14968 5040 15020
rect 6000 15036 6052 15088
rect 7380 15036 7432 15088
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 9220 15036 9272 15088
rect 10140 15079 10192 15088
rect 10140 15045 10149 15079
rect 10149 15045 10183 15079
rect 10183 15045 10192 15079
rect 10140 15036 10192 15045
rect 10600 15036 10652 15088
rect 12532 15079 12584 15088
rect 12532 15045 12541 15079
rect 12541 15045 12575 15079
rect 12575 15045 12584 15079
rect 12532 15036 12584 15045
rect 14924 15036 14976 15088
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 4620 14832 4672 14884
rect 7748 14968 7800 15020
rect 10692 15011 10744 15020
rect 6920 14900 6972 14952
rect 8208 14900 8260 14952
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 11520 14968 11572 15020
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12440 14968 12492 15020
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 14004 14968 14056 15020
rect 14280 14968 14332 15020
rect 12348 14943 12400 14952
rect 12348 14909 12374 14943
rect 12374 14909 12400 14943
rect 12348 14900 12400 14909
rect 12992 14900 13044 14952
rect 15660 14968 15712 15020
rect 17684 15036 17736 15088
rect 19708 15036 19760 15088
rect 16120 15011 16172 15020
rect 16120 14977 16129 15011
rect 16129 14977 16163 15011
rect 16163 14977 16172 15011
rect 16672 15011 16724 15020
rect 16120 14968 16172 14977
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 17500 14968 17552 15020
rect 17868 15011 17920 15020
rect 17868 14977 17877 15011
rect 17877 14977 17911 15011
rect 17911 14977 17920 15011
rect 17868 14968 17920 14977
rect 18236 14968 18288 15020
rect 16028 14900 16080 14952
rect 16856 14900 16908 14952
rect 19432 14968 19484 15020
rect 20352 15036 20404 15088
rect 8116 14832 8168 14884
rect 11980 14832 12032 14884
rect 16396 14832 16448 14884
rect 17776 14832 17828 14884
rect 18328 14832 18380 14884
rect 19248 14875 19300 14884
rect 19248 14841 19257 14875
rect 19257 14841 19291 14875
rect 19291 14841 19300 14875
rect 19248 14832 19300 14841
rect 2596 14764 2648 14816
rect 4804 14764 4856 14816
rect 5356 14764 5408 14816
rect 5724 14807 5776 14816
rect 5724 14773 5733 14807
rect 5733 14773 5767 14807
rect 5767 14773 5776 14807
rect 5724 14764 5776 14773
rect 6828 14764 6880 14816
rect 8392 14764 8444 14816
rect 8852 14764 8904 14816
rect 9680 14764 9732 14816
rect 10140 14764 10192 14816
rect 10416 14764 10468 14816
rect 13636 14764 13688 14816
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 17132 14764 17184 14816
rect 17592 14764 17644 14816
rect 20444 14764 20496 14816
rect 4338 14662 4390 14714
rect 4402 14662 4454 14714
rect 4466 14662 4518 14714
rect 4530 14662 4582 14714
rect 4594 14662 4646 14714
rect 11116 14662 11168 14714
rect 11180 14662 11232 14714
rect 11244 14662 11296 14714
rect 11308 14662 11360 14714
rect 11372 14662 11424 14714
rect 17893 14662 17945 14714
rect 17957 14662 18009 14714
rect 18021 14662 18073 14714
rect 18085 14662 18137 14714
rect 18149 14662 18201 14714
rect 3240 14560 3292 14612
rect 4252 14560 4304 14612
rect 2412 14492 2464 14544
rect 1768 14356 1820 14408
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2872 14399 2924 14408
rect 2596 14356 2648 14365
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 5080 14560 5132 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 6276 14560 6328 14612
rect 7564 14560 7616 14612
rect 9220 14560 9272 14612
rect 10048 14560 10100 14612
rect 12072 14560 12124 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14280 14560 14332 14612
rect 16856 14560 16908 14612
rect 17132 14603 17184 14612
rect 17132 14569 17141 14603
rect 17141 14569 17175 14603
rect 17175 14569 17184 14603
rect 17132 14560 17184 14569
rect 17776 14560 17828 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 20720 14603 20772 14612
rect 20720 14569 20729 14603
rect 20729 14569 20763 14603
rect 20763 14569 20772 14603
rect 20720 14560 20772 14569
rect 5172 14424 5224 14476
rect 7196 14467 7248 14476
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 5356 14356 5408 14408
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7380 14424 7432 14476
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 10784 14492 10836 14544
rect 10692 14467 10744 14476
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4988 14288 5040 14340
rect 5540 14288 5592 14340
rect 8852 14356 8904 14408
rect 9312 14356 9364 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 10692 14433 10701 14467
rect 10701 14433 10735 14467
rect 10735 14433 10744 14467
rect 10692 14424 10744 14433
rect 9864 14356 9916 14365
rect 10600 14399 10652 14408
rect 10600 14365 10609 14399
rect 10609 14365 10643 14399
rect 10643 14365 10652 14399
rect 10600 14356 10652 14365
rect 15476 14492 15528 14544
rect 12072 14424 12124 14476
rect 11980 14399 12032 14408
rect 11980 14365 11987 14399
rect 11987 14365 12032 14399
rect 11980 14356 12032 14365
rect 13452 14424 13504 14476
rect 13268 14399 13320 14408
rect 8852 14220 8904 14272
rect 9864 14220 9916 14272
rect 11704 14288 11756 14340
rect 12072 14331 12124 14340
rect 12072 14297 12081 14331
rect 12081 14297 12115 14331
rect 12115 14297 12124 14331
rect 12072 14288 12124 14297
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 13636 14356 13688 14408
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14740 14424 14792 14476
rect 19340 14424 19392 14476
rect 14372 14356 14424 14365
rect 16028 14356 16080 14408
rect 16120 14356 16172 14408
rect 16948 14356 17000 14408
rect 17500 14356 17552 14408
rect 18236 14356 18288 14408
rect 19616 14399 19668 14408
rect 10692 14220 10744 14272
rect 11796 14220 11848 14272
rect 14004 14288 14056 14340
rect 12256 14220 12308 14272
rect 13544 14220 13596 14272
rect 14280 14220 14332 14272
rect 14832 14220 14884 14272
rect 17132 14220 17184 14272
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20076 14356 20128 14408
rect 20536 14399 20588 14408
rect 18512 14288 18564 14340
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 20260 14288 20312 14340
rect 7727 14118 7779 14170
rect 7791 14118 7843 14170
rect 7855 14118 7907 14170
rect 7919 14118 7971 14170
rect 7983 14118 8035 14170
rect 14504 14118 14556 14170
rect 14568 14118 14620 14170
rect 14632 14118 14684 14170
rect 14696 14118 14748 14170
rect 14760 14118 14812 14170
rect 3332 14059 3384 14068
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 2964 13948 3016 14000
rect 3884 13948 3936 14000
rect 5356 14016 5408 14068
rect 6644 14016 6696 14068
rect 7656 14016 7708 14068
rect 8208 14016 8260 14068
rect 9956 14016 10008 14068
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 13452 14016 13504 14068
rect 16028 14016 16080 14068
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 17316 14016 17368 14068
rect 18236 14016 18288 14068
rect 19800 14016 19852 14068
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 20444 14016 20496 14068
rect 7196 13948 7248 14000
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 2780 13744 2832 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 2136 13719 2188 13728
rect 2136 13685 2145 13719
rect 2145 13685 2179 13719
rect 2179 13685 2188 13719
rect 2136 13676 2188 13685
rect 4160 13812 4212 13864
rect 3240 13744 3292 13796
rect 4988 13880 5040 13932
rect 5448 13880 5500 13932
rect 7472 13880 7524 13932
rect 8116 13991 8168 14000
rect 8116 13957 8125 13991
rect 8125 13957 8159 13991
rect 8159 13957 8168 13991
rect 8116 13948 8168 13957
rect 8852 13948 8904 14000
rect 11704 13948 11756 14000
rect 10140 13923 10192 13932
rect 5724 13812 5776 13864
rect 6828 13812 6880 13864
rect 5540 13744 5592 13796
rect 3700 13676 3752 13728
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 6920 13744 6972 13796
rect 8300 13812 8352 13864
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 10692 13923 10744 13932
rect 10692 13889 10701 13923
rect 10701 13889 10735 13923
rect 10735 13889 10744 13923
rect 10692 13880 10744 13889
rect 10416 13812 10468 13864
rect 10784 13812 10836 13864
rect 11980 13948 12032 14000
rect 12256 13948 12308 14000
rect 14188 13991 14240 14000
rect 14188 13957 14197 13991
rect 14197 13957 14231 13991
rect 14231 13957 14240 13991
rect 14188 13948 14240 13957
rect 12900 13880 12952 13932
rect 14004 13923 14056 13932
rect 8392 13744 8444 13796
rect 10968 13744 11020 13796
rect 11612 13744 11664 13796
rect 11980 13744 12032 13796
rect 12348 13744 12400 13796
rect 9036 13676 9088 13728
rect 9404 13676 9456 13728
rect 9588 13676 9640 13728
rect 9956 13676 10008 13728
rect 10784 13719 10836 13728
rect 10784 13685 10793 13719
rect 10793 13685 10827 13719
rect 10827 13685 10836 13719
rect 10784 13676 10836 13685
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 12072 13676 12124 13728
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 14832 13880 14884 13932
rect 18604 13948 18656 14000
rect 15200 13880 15252 13932
rect 15752 13880 15804 13932
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 17684 13880 17736 13932
rect 19248 13948 19300 14000
rect 19708 13948 19760 14000
rect 14004 13744 14056 13796
rect 18144 13855 18196 13864
rect 17684 13744 17736 13796
rect 18144 13821 18153 13855
rect 18153 13821 18187 13855
rect 18187 13821 18196 13855
rect 18144 13812 18196 13821
rect 18328 13812 18380 13864
rect 19340 13880 19392 13932
rect 19892 13880 19944 13932
rect 20168 13923 20220 13932
rect 20168 13889 20174 13923
rect 20174 13889 20208 13923
rect 20208 13889 20220 13923
rect 20168 13880 20220 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 20352 13812 20404 13864
rect 19524 13744 19576 13796
rect 18236 13676 18288 13728
rect 18512 13676 18564 13728
rect 19432 13676 19484 13728
rect 19800 13676 19852 13728
rect 4338 13574 4390 13626
rect 4402 13574 4454 13626
rect 4466 13574 4518 13626
rect 4530 13574 4582 13626
rect 4594 13574 4646 13626
rect 11116 13574 11168 13626
rect 11180 13574 11232 13626
rect 11244 13574 11296 13626
rect 11308 13574 11360 13626
rect 11372 13574 11424 13626
rect 17893 13574 17945 13626
rect 17957 13574 18009 13626
rect 18021 13574 18073 13626
rect 18085 13574 18137 13626
rect 18149 13574 18201 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 3148 13472 3200 13524
rect 3424 13472 3476 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 2136 13379 2188 13388
rect 2136 13345 2145 13379
rect 2145 13345 2179 13379
rect 2179 13345 2188 13379
rect 2136 13336 2188 13345
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 6460 13404 6512 13456
rect 7656 13404 7708 13456
rect 8576 13404 8628 13456
rect 9312 13472 9364 13524
rect 10048 13472 10100 13524
rect 2228 13336 2280 13345
rect 3332 13268 3384 13320
rect 3424 13268 3476 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 5080 13336 5132 13388
rect 5540 13336 5592 13388
rect 6644 13311 6696 13320
rect 2320 13132 2372 13184
rect 2688 13132 2740 13184
rect 4620 13132 4672 13184
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 5448 13200 5500 13252
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 7564 13336 7616 13388
rect 8116 13336 8168 13388
rect 8852 13336 8904 13388
rect 9128 13336 9180 13388
rect 9404 13404 9456 13456
rect 10140 13404 10192 13456
rect 10232 13404 10284 13456
rect 10048 13336 10100 13388
rect 10784 13404 10836 13456
rect 5816 13200 5868 13252
rect 7472 13268 7524 13320
rect 8392 13268 8444 13320
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 11796 13472 11848 13524
rect 12348 13472 12400 13524
rect 12900 13472 12952 13524
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 14924 13515 14976 13524
rect 14924 13481 14933 13515
rect 14933 13481 14967 13515
rect 14967 13481 14976 13515
rect 14924 13472 14976 13481
rect 17500 13472 17552 13524
rect 19708 13472 19760 13524
rect 20536 13472 20588 13524
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 18236 13404 18288 13456
rect 11244 13268 11296 13320
rect 12072 13268 12124 13320
rect 16120 13336 16172 13388
rect 16580 13379 16632 13388
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 7288 13200 7340 13252
rect 8852 13132 8904 13184
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 9220 13132 9272 13184
rect 11428 13200 11480 13252
rect 12348 13200 12400 13252
rect 14004 13200 14056 13252
rect 14280 13268 14332 13320
rect 14372 13200 14424 13252
rect 15476 13268 15528 13320
rect 15844 13200 15896 13252
rect 10232 13132 10284 13184
rect 10692 13132 10744 13184
rect 12624 13132 12676 13184
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 16580 13336 16632 13345
rect 16856 13336 16908 13388
rect 17132 13268 17184 13320
rect 17684 13200 17736 13252
rect 18052 13268 18104 13320
rect 20444 13404 20496 13456
rect 20628 13336 20680 13388
rect 19524 13268 19576 13320
rect 18512 13243 18564 13252
rect 18512 13209 18521 13243
rect 18521 13209 18555 13243
rect 18555 13209 18564 13243
rect 18512 13200 18564 13209
rect 18604 13200 18656 13252
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 16212 13132 16264 13184
rect 16856 13132 16908 13184
rect 18052 13132 18104 13184
rect 19432 13132 19484 13184
rect 20720 13200 20772 13252
rect 7727 13030 7779 13082
rect 7791 13030 7843 13082
rect 7855 13030 7907 13082
rect 7919 13030 7971 13082
rect 7983 13030 8035 13082
rect 14504 13030 14556 13082
rect 14568 13030 14620 13082
rect 14632 13030 14684 13082
rect 14696 13030 14748 13082
rect 14760 13030 14812 13082
rect 6552 12928 6604 12980
rect 2780 12860 2832 12912
rect 3792 12903 3844 12912
rect 3792 12869 3801 12903
rect 3801 12869 3835 12903
rect 3835 12869 3844 12903
rect 3792 12860 3844 12869
rect 5816 12860 5868 12912
rect 1860 12835 1912 12844
rect 1860 12801 1869 12835
rect 1869 12801 1903 12835
rect 1903 12801 1912 12835
rect 1860 12792 1912 12801
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 3240 12835 3292 12844
rect 2964 12792 3016 12801
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 4804 12792 4856 12844
rect 3148 12767 3200 12776
rect 3148 12733 3157 12767
rect 3157 12733 3191 12767
rect 3191 12733 3200 12767
rect 3148 12724 3200 12733
rect 3424 12724 3476 12776
rect 5172 12792 5224 12844
rect 5448 12792 5500 12844
rect 9772 12928 9824 12980
rect 10232 12971 10284 12980
rect 10232 12937 10241 12971
rect 10241 12937 10275 12971
rect 10275 12937 10284 12971
rect 10232 12928 10284 12937
rect 10416 12928 10468 12980
rect 7472 12903 7524 12912
rect 7472 12869 7481 12903
rect 7481 12869 7515 12903
rect 7515 12869 7524 12903
rect 7472 12860 7524 12869
rect 9128 12860 9180 12912
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 8852 12792 8904 12844
rect 9036 12792 9088 12844
rect 9588 12792 9640 12844
rect 10692 12860 10744 12912
rect 11704 12928 11756 12980
rect 14096 12928 14148 12980
rect 15016 12928 15068 12980
rect 17040 12928 17092 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 19984 12928 20036 12980
rect 11796 12860 11848 12912
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 5540 12724 5592 12776
rect 5632 12724 5684 12776
rect 6092 12724 6144 12776
rect 7472 12724 7524 12776
rect 14004 12792 14056 12844
rect 14188 12792 14240 12844
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 17408 12860 17460 12912
rect 20168 12860 20220 12912
rect 10692 12767 10744 12776
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 12808 12724 12860 12776
rect 13268 12724 13320 12776
rect 4620 12656 4672 12708
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6828 12588 6880 12640
rect 7196 12588 7248 12640
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 9128 12588 9180 12640
rect 9496 12656 9548 12708
rect 12624 12656 12676 12708
rect 15200 12724 15252 12776
rect 17316 12792 17368 12844
rect 17776 12792 17828 12844
rect 18328 12792 18380 12844
rect 19156 12792 19208 12844
rect 20352 12792 20404 12844
rect 17040 12724 17092 12776
rect 13544 12656 13596 12708
rect 16948 12656 17000 12708
rect 9864 12588 9916 12640
rect 10968 12588 11020 12640
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 13176 12588 13228 12640
rect 13912 12588 13964 12640
rect 14464 12588 14516 12640
rect 14740 12588 14792 12640
rect 17224 12588 17276 12640
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 20628 12631 20680 12640
rect 20628 12597 20637 12631
rect 20637 12597 20671 12631
rect 20671 12597 20680 12631
rect 20628 12588 20680 12597
rect 4338 12486 4390 12538
rect 4402 12486 4454 12538
rect 4466 12486 4518 12538
rect 4530 12486 4582 12538
rect 4594 12486 4646 12538
rect 11116 12486 11168 12538
rect 11180 12486 11232 12538
rect 11244 12486 11296 12538
rect 11308 12486 11360 12538
rect 11372 12486 11424 12538
rect 17893 12486 17945 12538
rect 17957 12486 18009 12538
rect 18021 12486 18073 12538
rect 18085 12486 18137 12538
rect 18149 12486 18201 12538
rect 1492 12384 1544 12436
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 5540 12384 5592 12436
rect 7288 12384 7340 12436
rect 3792 12316 3844 12368
rect 6184 12359 6236 12368
rect 6184 12325 6193 12359
rect 6193 12325 6227 12359
rect 6227 12325 6236 12359
rect 6184 12316 6236 12325
rect 3056 12248 3108 12300
rect 3240 12291 3292 12300
rect 3240 12257 3249 12291
rect 3249 12257 3283 12291
rect 3283 12257 3292 12291
rect 3240 12248 3292 12257
rect 4896 12248 4948 12300
rect 5264 12291 5316 12300
rect 5264 12257 5273 12291
rect 5273 12257 5307 12291
rect 5307 12257 5316 12291
rect 5264 12248 5316 12257
rect 5356 12248 5408 12300
rect 1400 12180 1452 12232
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 6000 12223 6052 12232
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 6000 12180 6052 12189
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 6828 12180 6880 12232
rect 7196 12180 7248 12232
rect 7564 12180 7616 12232
rect 9496 12384 9548 12436
rect 11980 12384 12032 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 13452 12427 13504 12436
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 14004 12384 14056 12436
rect 8208 12316 8260 12368
rect 15016 12384 15068 12436
rect 15200 12384 15252 12436
rect 16028 12384 16080 12436
rect 16580 12384 16632 12436
rect 17316 12384 17368 12436
rect 17684 12384 17736 12436
rect 19800 12384 19852 12436
rect 19984 12384 20036 12436
rect 8116 12248 8168 12300
rect 12900 12248 12952 12300
rect 14188 12248 14240 12300
rect 2964 12112 3016 12164
rect 10692 12180 10744 12232
rect 10784 12223 10836 12232
rect 10784 12189 10818 12223
rect 10818 12189 10836 12223
rect 10784 12180 10836 12189
rect 11612 12180 11664 12232
rect 12072 12180 12124 12232
rect 13544 12180 13596 12232
rect 13912 12180 13964 12232
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 15936 12316 15988 12368
rect 14556 12291 14608 12300
rect 14556 12257 14565 12291
rect 14565 12257 14599 12291
rect 14599 12257 14608 12291
rect 14556 12248 14608 12257
rect 15660 12248 15712 12300
rect 13084 12112 13136 12164
rect 2596 12044 2648 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 4068 12044 4120 12096
rect 5356 12044 5408 12096
rect 8300 12044 8352 12096
rect 10876 12044 10928 12096
rect 14740 12180 14792 12232
rect 14832 12180 14884 12232
rect 15752 12112 15804 12164
rect 19524 12316 19576 12368
rect 20628 12248 20680 12300
rect 16212 12180 16264 12232
rect 16856 12180 16908 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17684 12223 17736 12232
rect 17408 12180 17460 12189
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 17868 12180 17920 12232
rect 19708 12180 19760 12232
rect 20352 12180 20404 12232
rect 19892 12112 19944 12164
rect 17500 12044 17552 12096
rect 18144 12044 18196 12096
rect 19248 12044 19300 12096
rect 7727 11942 7779 11994
rect 7791 11942 7843 11994
rect 7855 11942 7907 11994
rect 7919 11942 7971 11994
rect 7983 11942 8035 11994
rect 14504 11942 14556 11994
rect 14568 11942 14620 11994
rect 14632 11942 14684 11994
rect 14696 11942 14748 11994
rect 14760 11942 14812 11994
rect 2136 11840 2188 11892
rect 2688 11840 2740 11892
rect 5356 11883 5408 11892
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 2872 11704 2924 11756
rect 3884 11772 3936 11824
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 8668 11840 8720 11892
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 12532 11840 12584 11892
rect 15200 11840 15252 11892
rect 15292 11840 15344 11892
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 19156 11840 19208 11892
rect 19524 11840 19576 11892
rect 7104 11772 7156 11824
rect 3976 11704 4028 11756
rect 4068 11704 4120 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 4804 11636 4856 11688
rect 5356 11636 5408 11688
rect 6184 11636 6236 11688
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 9772 11772 9824 11824
rect 10140 11772 10192 11824
rect 9312 11704 9364 11756
rect 10416 11679 10468 11688
rect 10416 11645 10425 11679
rect 10425 11645 10459 11679
rect 10459 11645 10468 11679
rect 10416 11636 10468 11645
rect 9128 11568 9180 11620
rect 10876 11704 10928 11756
rect 12072 11704 12124 11756
rect 10968 11636 11020 11688
rect 12716 11704 12768 11756
rect 15108 11772 15160 11824
rect 18144 11772 18196 11824
rect 18972 11772 19024 11824
rect 14648 11747 14700 11756
rect 12900 11636 12952 11688
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 14832 11704 14884 11756
rect 15384 11704 15436 11756
rect 12256 11568 12308 11620
rect 15292 11636 15344 11688
rect 13636 11568 13688 11620
rect 16304 11704 16356 11756
rect 17684 11704 17736 11756
rect 17776 11704 17828 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18512 11704 18564 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 20168 11772 20220 11824
rect 20536 11772 20588 11824
rect 18604 11704 18656 11713
rect 18144 11636 18196 11688
rect 20260 11636 20312 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2872 11500 2924 11552
rect 4160 11500 4212 11552
rect 4252 11500 4304 11552
rect 7656 11500 7708 11552
rect 8944 11500 8996 11552
rect 9588 11500 9640 11552
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12992 11543 13044 11552
rect 12440 11500 12492 11509
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 13084 11500 13136 11552
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 14556 11500 14608 11552
rect 16856 11568 16908 11620
rect 17408 11568 17460 11620
rect 17684 11568 17736 11620
rect 17868 11568 17920 11620
rect 18696 11568 18748 11620
rect 15660 11500 15712 11552
rect 17592 11500 17644 11552
rect 19524 11543 19576 11552
rect 19524 11509 19533 11543
rect 19533 11509 19567 11543
rect 19567 11509 19576 11543
rect 19524 11500 19576 11509
rect 4338 11398 4390 11450
rect 4402 11398 4454 11450
rect 4466 11398 4518 11450
rect 4530 11398 4582 11450
rect 4594 11398 4646 11450
rect 11116 11398 11168 11450
rect 11180 11398 11232 11450
rect 11244 11398 11296 11450
rect 11308 11398 11360 11450
rect 11372 11398 11424 11450
rect 17893 11398 17945 11450
rect 17957 11398 18009 11450
rect 18021 11398 18073 11450
rect 18085 11398 18137 11450
rect 18149 11398 18201 11450
rect 2688 11296 2740 11348
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 4712 11296 4764 11348
rect 6276 11296 6328 11348
rect 7196 11339 7248 11348
rect 7196 11305 7205 11339
rect 7205 11305 7239 11339
rect 7239 11305 7248 11339
rect 7196 11296 7248 11305
rect 9312 11296 9364 11348
rect 10324 11339 10376 11348
rect 3700 11228 3752 11280
rect 6920 11228 6972 11280
rect 8760 11228 8812 11280
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 10692 11296 10744 11348
rect 10968 11296 11020 11348
rect 11520 11296 11572 11348
rect 12072 11296 12124 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 12992 11296 13044 11348
rect 13452 11296 13504 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 15476 11296 15528 11348
rect 17776 11296 17828 11348
rect 2872 11160 2924 11212
rect 2412 11092 2464 11144
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 2688 11092 2740 11144
rect 2780 11092 2832 11144
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 2228 11024 2280 11076
rect 3332 11024 3384 11076
rect 4712 11160 4764 11212
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 5632 11092 5684 11144
rect 5816 11092 5868 11144
rect 5724 11024 5776 11076
rect 7196 11092 7248 11144
rect 7656 11092 7708 11144
rect 6276 11024 6328 11076
rect 9128 11092 9180 11144
rect 9772 11092 9824 11144
rect 10784 11092 10836 11144
rect 12348 11092 12400 11144
rect 14648 11228 14700 11280
rect 12900 11160 12952 11212
rect 14096 11160 14148 11212
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13636 11092 13688 11144
rect 15292 11160 15344 11212
rect 16028 11228 16080 11280
rect 16856 11228 16908 11280
rect 15844 11160 15896 11212
rect 17592 11203 17644 11212
rect 8576 11024 8628 11076
rect 9588 11024 9640 11076
rect 12440 11024 12492 11076
rect 14556 11024 14608 11076
rect 16304 11092 16356 11144
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 14832 11024 14884 11076
rect 16764 11092 16816 11144
rect 17132 11092 17184 11144
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 18972 11092 19024 11144
rect 19340 11160 19392 11212
rect 19800 11160 19852 11212
rect 19432 11092 19484 11144
rect 2688 10999 2740 11008
rect 2688 10965 2697 10999
rect 2697 10965 2731 10999
rect 2731 10965 2740 10999
rect 2688 10956 2740 10965
rect 6920 10956 6972 11008
rect 8208 10956 8260 11008
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 12256 10956 12308 11008
rect 15200 10956 15252 11008
rect 15660 10956 15712 11008
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 16396 10956 16448 11008
rect 17592 11024 17644 11076
rect 18696 11067 18748 11076
rect 18696 11033 18705 11067
rect 18705 11033 18739 11067
rect 18739 11033 18748 11067
rect 18696 11024 18748 11033
rect 19340 10956 19392 11008
rect 19984 10999 20036 11008
rect 19984 10965 19993 10999
rect 19993 10965 20027 10999
rect 20027 10965 20036 10999
rect 19984 10956 20036 10965
rect 20076 10999 20128 11008
rect 20076 10965 20085 10999
rect 20085 10965 20119 10999
rect 20119 10965 20128 10999
rect 20076 10956 20128 10965
rect 7727 10854 7779 10906
rect 7791 10854 7843 10906
rect 7855 10854 7907 10906
rect 7919 10854 7971 10906
rect 7983 10854 8035 10906
rect 14504 10854 14556 10906
rect 14568 10854 14620 10906
rect 14632 10854 14684 10906
rect 14696 10854 14748 10906
rect 14760 10854 14812 10906
rect 2044 10752 2096 10804
rect 2504 10752 2556 10804
rect 2228 10684 2280 10736
rect 2780 10684 2832 10736
rect 3976 10752 4028 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3332 10616 3384 10668
rect 4804 10752 4856 10804
rect 5632 10752 5684 10804
rect 7656 10752 7708 10804
rect 8668 10752 8720 10804
rect 14832 10752 14884 10804
rect 16304 10752 16356 10804
rect 18512 10795 18564 10804
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 19984 10752 20036 10804
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 4160 10616 4212 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 5632 10659 5684 10668
rect 4252 10548 4304 10600
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 8944 10684 8996 10736
rect 12808 10727 12860 10736
rect 12808 10693 12817 10727
rect 12817 10693 12851 10727
rect 12851 10693 12860 10727
rect 12808 10684 12860 10693
rect 13544 10684 13596 10736
rect 6828 10548 6880 10600
rect 7656 10616 7708 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 8208 10616 8260 10668
rect 10048 10659 10100 10668
rect 9220 10548 9272 10600
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10692 10616 10744 10668
rect 12992 10616 13044 10668
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 16120 10684 16172 10736
rect 18604 10684 18656 10736
rect 14648 10616 14700 10668
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 17776 10616 17828 10668
rect 19340 10684 19392 10736
rect 19064 10659 19116 10668
rect 10876 10548 10928 10600
rect 11704 10548 11756 10600
rect 13636 10548 13688 10600
rect 8944 10480 8996 10532
rect 9864 10480 9916 10532
rect 10416 10480 10468 10532
rect 13728 10480 13780 10532
rect 14188 10480 14240 10532
rect 17684 10548 17736 10600
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 19616 10616 19668 10668
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 19524 10548 19576 10600
rect 19984 10548 20036 10600
rect 20628 10548 20680 10600
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2964 10412 3016 10464
rect 6644 10412 6696 10464
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 7564 10455 7616 10464
rect 6828 10412 6880 10421
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 7656 10412 7708 10464
rect 8116 10412 8168 10464
rect 8668 10412 8720 10464
rect 9220 10412 9272 10464
rect 10600 10412 10652 10464
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 15844 10412 15896 10464
rect 16488 10412 16540 10464
rect 17224 10412 17276 10464
rect 19616 10412 19668 10464
rect 19892 10412 19944 10464
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 4338 10310 4390 10362
rect 4402 10310 4454 10362
rect 4466 10310 4518 10362
rect 4530 10310 4582 10362
rect 4594 10310 4646 10362
rect 11116 10310 11168 10362
rect 11180 10310 11232 10362
rect 11244 10310 11296 10362
rect 11308 10310 11360 10362
rect 11372 10310 11424 10362
rect 17893 10310 17945 10362
rect 17957 10310 18009 10362
rect 18021 10310 18073 10362
rect 18085 10310 18137 10362
rect 18149 10310 18201 10362
rect 2504 10208 2556 10260
rect 4160 10208 4212 10260
rect 7288 10208 7340 10260
rect 7840 10208 7892 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8944 10251 8996 10260
rect 8300 10208 8352 10217
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 6460 10140 6512 10192
rect 6920 10072 6972 10124
rect 9404 10208 9456 10260
rect 9496 10208 9548 10260
rect 10048 10208 10100 10260
rect 10416 10208 10468 10260
rect 12348 10208 12400 10260
rect 12624 10208 12676 10260
rect 13268 10208 13320 10260
rect 13728 10208 13780 10260
rect 12992 10140 13044 10192
rect 14556 10208 14608 10260
rect 16488 10140 16540 10192
rect 19524 10208 19576 10260
rect 19892 10208 19944 10260
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 19984 10183 20036 10192
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 16672 10072 16724 10124
rect 2412 10004 2464 10056
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2872 10047 2924 10056
rect 2596 10004 2648 10013
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3884 10047 3936 10056
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 5080 10004 5132 10056
rect 5448 10004 5500 10056
rect 5632 10004 5684 10056
rect 7564 10004 7616 10056
rect 8116 10004 8168 10056
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 11428 10004 11480 10056
rect 12532 10004 12584 10056
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 6276 9868 6328 9920
rect 8944 9868 8996 9920
rect 9496 9868 9548 9920
rect 10140 9868 10192 9920
rect 11612 9936 11664 9988
rect 13820 10004 13872 10056
rect 19984 10149 19993 10183
rect 19993 10149 20027 10183
rect 20027 10149 20036 10183
rect 19984 10140 20036 10149
rect 14372 9936 14424 9988
rect 14648 9979 14700 9988
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 15016 9936 15068 9988
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 13084 9868 13136 9920
rect 13728 9868 13780 9920
rect 14004 9868 14056 9920
rect 16212 9936 16264 9988
rect 16672 9936 16724 9988
rect 17224 9936 17276 9988
rect 17500 9979 17552 9988
rect 17500 9945 17509 9979
rect 17509 9945 17543 9979
rect 17543 9945 17552 9979
rect 20260 10072 20312 10124
rect 19340 10004 19392 10056
rect 20628 10004 20680 10056
rect 17500 9936 17552 9945
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 7727 9766 7779 9818
rect 7791 9766 7843 9818
rect 7855 9766 7907 9818
rect 7919 9766 7971 9818
rect 7983 9766 8035 9818
rect 14504 9766 14556 9818
rect 14568 9766 14620 9818
rect 14632 9766 14684 9818
rect 14696 9766 14748 9818
rect 14760 9766 14812 9818
rect 1400 9528 1452 9580
rect 2964 9596 3016 9648
rect 5448 9664 5500 9716
rect 6368 9664 6420 9716
rect 6828 9664 6880 9716
rect 6920 9664 6972 9716
rect 7104 9596 7156 9648
rect 8300 9664 8352 9716
rect 9496 9664 9548 9716
rect 10048 9664 10100 9716
rect 13820 9664 13872 9716
rect 14280 9664 14332 9716
rect 17500 9664 17552 9716
rect 2688 9528 2740 9580
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3424 9528 3476 9580
rect 1768 9460 1820 9512
rect 1860 9460 1912 9512
rect 1492 9435 1544 9444
rect 1492 9401 1501 9435
rect 1501 9401 1535 9435
rect 1535 9401 1544 9435
rect 1492 9392 1544 9401
rect 5356 9528 5408 9580
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 6092 9528 6144 9580
rect 7012 9528 7064 9580
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 8576 9596 8628 9648
rect 12348 9596 12400 9648
rect 8668 9528 8720 9580
rect 11428 9528 11480 9580
rect 12256 9528 12308 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 14004 9528 14056 9580
rect 14372 9596 14424 9648
rect 17408 9596 17460 9648
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 7380 9460 7432 9512
rect 9036 9460 9088 9512
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4988 9324 5040 9376
rect 6000 9392 6052 9444
rect 8300 9392 8352 9444
rect 9588 9392 9640 9444
rect 11980 9460 12032 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 13728 9460 13780 9512
rect 17500 9528 17552 9580
rect 18052 9528 18104 9580
rect 18604 9596 18656 9648
rect 18696 9596 18748 9648
rect 18512 9528 18564 9580
rect 19248 9460 19300 9512
rect 11796 9392 11848 9444
rect 5632 9324 5684 9376
rect 6184 9324 6236 9376
rect 6828 9324 6880 9376
rect 10416 9324 10468 9376
rect 10600 9324 10652 9376
rect 12624 9324 12676 9376
rect 12716 9324 12768 9376
rect 17224 9392 17276 9444
rect 19800 9392 19852 9444
rect 14832 9324 14884 9376
rect 16304 9324 16356 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 19708 9367 19760 9376
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 4338 9222 4390 9274
rect 4402 9222 4454 9274
rect 4466 9222 4518 9274
rect 4530 9222 4582 9274
rect 4594 9222 4646 9274
rect 11116 9222 11168 9274
rect 11180 9222 11232 9274
rect 11244 9222 11296 9274
rect 11308 9222 11360 9274
rect 11372 9222 11424 9274
rect 17893 9222 17945 9274
rect 17957 9222 18009 9274
rect 18021 9222 18073 9274
rect 18085 9222 18137 9274
rect 18149 9222 18201 9274
rect 6092 9120 6144 9172
rect 8944 9120 8996 9172
rect 9496 9120 9548 9172
rect 10876 9120 10928 9172
rect 14372 9120 14424 9172
rect 15108 9120 15160 9172
rect 17500 9120 17552 9172
rect 18512 9120 18564 9172
rect 7380 9095 7432 9104
rect 7380 9061 7389 9095
rect 7389 9061 7423 9095
rect 7423 9061 7432 9095
rect 7380 9052 7432 9061
rect 10416 9052 10468 9104
rect 15384 9052 15436 9104
rect 16672 9052 16724 9104
rect 18696 9052 18748 9104
rect 3700 8984 3752 9036
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5172 9027 5224 9036
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 5264 8984 5316 9036
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 7104 8984 7156 9036
rect 7656 8984 7708 9036
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 3148 8916 3200 8968
rect 4160 8916 4212 8968
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6736 8916 6788 8968
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 6000 8848 6052 8900
rect 6920 8848 6972 8900
rect 7472 8848 7524 8900
rect 7748 8916 7800 8968
rect 10692 8984 10744 9036
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 11704 8984 11756 9036
rect 12256 8984 12308 9036
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 12532 8916 12584 8968
rect 12716 8916 12768 8968
rect 16764 8984 16816 9036
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 19892 9027 19944 9036
rect 18144 8984 18196 8993
rect 14372 8916 14424 8968
rect 10324 8848 10376 8900
rect 15844 8916 15896 8968
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 3608 8780 3660 8832
rect 3792 8780 3844 8832
rect 3976 8780 4028 8832
rect 5356 8780 5408 8832
rect 8116 8780 8168 8832
rect 10876 8780 10928 8832
rect 13268 8780 13320 8832
rect 14096 8780 14148 8832
rect 15292 8780 15344 8832
rect 16028 8848 16080 8900
rect 16488 8916 16540 8968
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 18236 8916 18288 8968
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 19708 8916 19760 8968
rect 20720 8891 20772 8900
rect 20720 8857 20729 8891
rect 20729 8857 20763 8891
rect 20763 8857 20772 8891
rect 20720 8848 20772 8857
rect 17500 8780 17552 8832
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 19524 8780 19576 8832
rect 19800 8780 19852 8832
rect 7727 8678 7779 8730
rect 7791 8678 7843 8730
rect 7855 8678 7907 8730
rect 7919 8678 7971 8730
rect 7983 8678 8035 8730
rect 14504 8678 14556 8730
rect 14568 8678 14620 8730
rect 14632 8678 14684 8730
rect 14696 8678 14748 8730
rect 14760 8678 14812 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 2504 8576 2556 8628
rect 2872 8551 2924 8560
rect 2872 8517 2881 8551
rect 2881 8517 2915 8551
rect 2915 8517 2924 8551
rect 2872 8508 2924 8517
rect 3792 8508 3844 8560
rect 2780 8440 2832 8492
rect 2504 8372 2556 8424
rect 3884 8440 3936 8492
rect 4712 8576 4764 8628
rect 5356 8619 5408 8628
rect 4252 8508 4304 8560
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 6736 8619 6788 8628
rect 6736 8585 6745 8619
rect 6745 8585 6779 8619
rect 6779 8585 6788 8619
rect 6736 8576 6788 8585
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 5540 8508 5592 8560
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 3148 8372 3200 8424
rect 4988 8440 5040 8492
rect 7656 8508 7708 8560
rect 7472 8483 7524 8492
rect 5172 8372 5224 8424
rect 6368 8372 6420 8424
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 4068 8304 4120 8356
rect 8116 8372 8168 8424
rect 1952 8279 2004 8288
rect 1952 8245 1961 8279
rect 1961 8245 1995 8279
rect 1995 8245 2004 8279
rect 1952 8236 2004 8245
rect 3792 8236 3844 8288
rect 6644 8236 6696 8288
rect 7472 8304 7524 8356
rect 9496 8508 9548 8560
rect 9956 8551 10008 8560
rect 8760 8440 8812 8492
rect 9956 8517 9965 8551
rect 9965 8517 9999 8551
rect 9999 8517 10008 8551
rect 9956 8508 10008 8517
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 13912 8576 13964 8628
rect 14004 8576 14056 8628
rect 15108 8576 15160 8628
rect 17960 8576 18012 8628
rect 19156 8576 19208 8628
rect 14832 8508 14884 8560
rect 14924 8508 14976 8560
rect 16396 8508 16448 8560
rect 16856 8508 16908 8560
rect 10784 8483 10836 8492
rect 10048 8304 10100 8356
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 13728 8440 13780 8492
rect 14188 8440 14240 8492
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11796 8372 11848 8424
rect 12808 8372 12860 8424
rect 15108 8440 15160 8492
rect 15476 8483 15528 8492
rect 15200 8372 15252 8424
rect 14832 8304 14884 8356
rect 15108 8347 15160 8356
rect 15108 8313 15117 8347
rect 15117 8313 15151 8347
rect 15151 8313 15160 8347
rect 15108 8304 15160 8313
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 15660 8372 15712 8424
rect 16120 8440 16172 8492
rect 16488 8440 16540 8492
rect 18328 8440 18380 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 15844 8372 15896 8424
rect 17592 8372 17644 8424
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 17040 8304 17092 8356
rect 17132 8304 17184 8356
rect 18604 8304 18656 8356
rect 9312 8236 9364 8288
rect 11704 8236 11756 8288
rect 13360 8236 13412 8288
rect 14924 8236 14976 8288
rect 16672 8236 16724 8288
rect 19156 8236 19208 8288
rect 4338 8134 4390 8186
rect 4402 8134 4454 8186
rect 4466 8134 4518 8186
rect 4530 8134 4582 8186
rect 4594 8134 4646 8186
rect 11116 8134 11168 8186
rect 11180 8134 11232 8186
rect 11244 8134 11296 8186
rect 11308 8134 11360 8186
rect 11372 8134 11424 8186
rect 17893 8134 17945 8186
rect 17957 8134 18009 8186
rect 18021 8134 18073 8186
rect 18085 8134 18137 8186
rect 18149 8134 18201 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 9128 8032 9180 8084
rect 9956 8032 10008 8084
rect 4988 7964 5040 8016
rect 5448 8007 5500 8016
rect 5448 7973 5457 8007
rect 5457 7973 5491 8007
rect 5491 7973 5500 8007
rect 5448 7964 5500 7973
rect 9772 8007 9824 8016
rect 2136 7896 2188 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 4160 7896 4212 7948
rect 3884 7828 3936 7880
rect 3976 7828 4028 7880
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5264 7828 5316 7880
rect 1952 7760 2004 7812
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 3700 7692 3752 7744
rect 5448 7692 5500 7744
rect 6736 7896 6788 7948
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 9772 7973 9781 8007
rect 9781 7973 9815 8007
rect 9815 7973 9824 8007
rect 9772 7964 9824 7973
rect 10140 7964 10192 8016
rect 7840 7896 7892 7905
rect 7380 7828 7432 7880
rect 10232 7896 10284 7948
rect 8576 7828 8628 7880
rect 9036 7828 9088 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 9680 7828 9732 7880
rect 10324 7828 10376 7880
rect 11704 7896 11756 7948
rect 10876 7828 10928 7880
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 12440 8032 12492 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 15476 8032 15528 8084
rect 15660 8032 15712 8084
rect 16672 8032 16724 8084
rect 16764 8032 16816 8084
rect 12808 7964 12860 8016
rect 15936 7964 15988 8016
rect 16120 7964 16172 8016
rect 19432 8032 19484 8084
rect 20260 8032 20312 8084
rect 17500 7964 17552 8016
rect 18328 7964 18380 8016
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12256 7828 12308 7880
rect 8852 7760 8904 7812
rect 6184 7692 6236 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 10508 7692 10560 7744
rect 11152 7692 11204 7744
rect 11704 7760 11756 7812
rect 12624 7828 12676 7880
rect 12808 7828 12860 7880
rect 13268 7828 13320 7880
rect 12532 7760 12584 7812
rect 13912 7828 13964 7880
rect 15016 7828 15068 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 13728 7692 13780 7744
rect 16304 7896 16356 7948
rect 16764 7896 16816 7948
rect 17868 7896 17920 7948
rect 19524 7964 19576 8016
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 17040 7828 17092 7880
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 18236 7828 18288 7880
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18788 7828 18840 7880
rect 19064 7828 19116 7880
rect 16672 7760 16724 7812
rect 20536 7803 20588 7812
rect 15476 7692 15528 7744
rect 15752 7692 15804 7744
rect 17960 7692 18012 7744
rect 18512 7692 18564 7744
rect 18604 7692 18656 7744
rect 18972 7692 19024 7744
rect 19340 7692 19392 7744
rect 20536 7769 20545 7803
rect 20545 7769 20579 7803
rect 20579 7769 20588 7803
rect 20536 7760 20588 7769
rect 20628 7735 20680 7744
rect 20628 7701 20637 7735
rect 20637 7701 20671 7735
rect 20671 7701 20680 7735
rect 20628 7692 20680 7701
rect 7727 7590 7779 7642
rect 7791 7590 7843 7642
rect 7855 7590 7907 7642
rect 7919 7590 7971 7642
rect 7983 7590 8035 7642
rect 14504 7590 14556 7642
rect 14568 7590 14620 7642
rect 14632 7590 14684 7642
rect 14696 7590 14748 7642
rect 14760 7590 14812 7642
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 6736 7488 6788 7540
rect 7472 7488 7524 7540
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 3792 7352 3844 7404
rect 5264 7420 5316 7472
rect 6552 7420 6604 7472
rect 9588 7488 9640 7540
rect 10140 7488 10192 7540
rect 10692 7488 10744 7540
rect 12256 7488 12308 7540
rect 13636 7531 13688 7540
rect 4252 7352 4304 7404
rect 4712 7352 4764 7404
rect 5356 7352 5408 7404
rect 5908 7352 5960 7404
rect 6368 7352 6420 7404
rect 10784 7420 10836 7472
rect 8300 7395 8352 7404
rect 3884 7216 3936 7268
rect 4896 7284 4948 7336
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8760 7352 8812 7404
rect 9588 7352 9640 7404
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 10600 7352 10652 7404
rect 11244 7352 11296 7404
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 9680 7284 9732 7336
rect 4160 7216 4212 7268
rect 10416 7284 10468 7336
rect 10232 7216 10284 7268
rect 11980 7352 12032 7404
rect 12256 7352 12308 7404
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 17868 7488 17920 7540
rect 18328 7488 18380 7540
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13820 7352 13872 7404
rect 13912 7352 13964 7404
rect 14924 7395 14976 7404
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15476 7352 15528 7404
rect 15108 7284 15160 7336
rect 15200 7284 15252 7336
rect 16028 7352 16080 7404
rect 16488 7352 16540 7404
rect 19064 7463 19116 7472
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17132 7352 17184 7404
rect 18144 7352 18196 7404
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 19064 7429 19073 7463
rect 19073 7429 19107 7463
rect 19107 7429 19116 7463
rect 19064 7420 19116 7429
rect 18604 7352 18656 7404
rect 18880 7352 18932 7404
rect 19156 7352 19208 7404
rect 3976 7148 4028 7200
rect 6000 7148 6052 7200
rect 6736 7191 6788 7200
rect 6736 7157 6745 7191
rect 6745 7157 6779 7191
rect 6779 7157 6788 7191
rect 6736 7148 6788 7157
rect 7196 7148 7248 7200
rect 9312 7148 9364 7200
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 13544 7216 13596 7268
rect 15384 7216 15436 7268
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13728 7148 13780 7200
rect 15292 7148 15344 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 15752 7148 15804 7200
rect 16304 7148 16356 7200
rect 20168 7284 20220 7336
rect 20260 7216 20312 7268
rect 18604 7148 18656 7200
rect 19892 7148 19944 7200
rect 4338 7046 4390 7098
rect 4402 7046 4454 7098
rect 4466 7046 4518 7098
rect 4530 7046 4582 7098
rect 4594 7046 4646 7098
rect 11116 7046 11168 7098
rect 11180 7046 11232 7098
rect 11244 7046 11296 7098
rect 11308 7046 11360 7098
rect 11372 7046 11424 7098
rect 17893 7046 17945 7098
rect 17957 7046 18009 7098
rect 18021 7046 18073 7098
rect 18085 7046 18137 7098
rect 18149 7046 18201 7098
rect 2872 6987 2924 6996
rect 2872 6953 2881 6987
rect 2881 6953 2915 6987
rect 2915 6953 2924 6987
rect 2872 6944 2924 6953
rect 3792 6944 3844 6996
rect 4252 6944 4304 6996
rect 5356 6944 5408 6996
rect 3516 6808 3568 6860
rect 2320 6740 2372 6792
rect 4252 6808 4304 6860
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3976 6740 4028 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 8300 6944 8352 6996
rect 10140 6944 10192 6996
rect 10692 6944 10744 6996
rect 12164 6944 12216 6996
rect 16028 6987 16080 6996
rect 6920 6876 6972 6928
rect 7288 6876 7340 6928
rect 7104 6808 7156 6860
rect 7656 6808 7708 6860
rect 8116 6876 8168 6928
rect 14372 6876 14424 6928
rect 16028 6953 16037 6987
rect 16037 6953 16071 6987
rect 16071 6953 16080 6987
rect 16028 6944 16080 6953
rect 16488 6944 16540 6996
rect 18420 6944 18472 6996
rect 18788 6944 18840 6996
rect 20168 6987 20220 6996
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7380 6740 7432 6792
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 9588 6808 9640 6860
rect 10416 6808 10468 6860
rect 11612 6808 11664 6860
rect 11980 6808 12032 6860
rect 15660 6876 15712 6928
rect 18696 6876 18748 6928
rect 19156 6876 19208 6928
rect 15016 6808 15068 6860
rect 17040 6808 17092 6860
rect 19340 6808 19392 6860
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9220 6740 9272 6792
rect 10968 6783 11020 6792
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 2596 6604 2648 6656
rect 8392 6672 8444 6724
rect 9588 6715 9640 6724
rect 4160 6604 4212 6656
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 5540 6604 5592 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9588 6681 9597 6715
rect 9597 6681 9631 6715
rect 9631 6681 9640 6715
rect 9588 6672 9640 6681
rect 9864 6672 9916 6724
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 11704 6740 11756 6792
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 13268 6783 13320 6792
rect 9956 6647 10008 6656
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11612 6672 11664 6724
rect 12164 6672 12216 6724
rect 12440 6672 12492 6724
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13728 6740 13780 6792
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 15660 6740 15712 6792
rect 15752 6740 15804 6792
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 16856 6740 16908 6792
rect 13452 6672 13504 6724
rect 14832 6672 14884 6724
rect 12716 6604 12768 6656
rect 14372 6604 14424 6656
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18696 6783 18748 6792
rect 18420 6740 18472 6749
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 19064 6740 19116 6792
rect 20076 6783 20128 6792
rect 19156 6672 19208 6724
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 15016 6604 15068 6613
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 17960 6604 18012 6656
rect 18328 6604 18380 6656
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 20628 6604 20680 6656
rect 7727 6502 7779 6554
rect 7791 6502 7843 6554
rect 7855 6502 7907 6554
rect 7919 6502 7971 6554
rect 7983 6502 8035 6554
rect 14504 6502 14556 6554
rect 14568 6502 14620 6554
rect 14632 6502 14684 6554
rect 14696 6502 14748 6554
rect 14760 6502 14812 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 3148 6400 3200 6452
rect 5172 6400 5224 6452
rect 6460 6400 6512 6452
rect 7380 6400 7432 6452
rect 9496 6443 9548 6452
rect 2504 6332 2556 6384
rect 1768 6264 1820 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2596 6307 2648 6316
rect 2320 6264 2372 6273
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 2964 6264 3016 6316
rect 4620 6332 4672 6384
rect 2872 6196 2924 6248
rect 3792 6264 3844 6316
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4712 6264 4764 6316
rect 4896 6264 4948 6316
rect 4988 6264 5040 6316
rect 7196 6264 7248 6316
rect 2964 6128 3016 6180
rect 4804 6196 4856 6248
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 10876 6443 10928 6452
rect 10876 6409 10885 6443
rect 10885 6409 10919 6443
rect 10919 6409 10928 6443
rect 10876 6400 10928 6409
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 10600 6332 10652 6384
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 9036 6307 9088 6316
rect 8392 6264 8444 6273
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 6920 6196 6972 6205
rect 10692 6264 10744 6316
rect 11612 6264 11664 6316
rect 6092 6128 6144 6180
rect 10968 6196 11020 6248
rect 12164 6400 12216 6452
rect 15016 6400 15068 6452
rect 12348 6332 12400 6384
rect 13268 6332 13320 6384
rect 14648 6332 14700 6384
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 14280 6264 14332 6316
rect 2136 6060 2188 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4160 6060 4212 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 6276 6060 6328 6112
rect 6736 6060 6788 6112
rect 6920 6060 6972 6112
rect 7380 6060 7432 6112
rect 8300 6060 8352 6112
rect 10600 6128 10652 6180
rect 10784 6060 10836 6112
rect 10968 6060 11020 6112
rect 13268 6196 13320 6248
rect 14924 6264 14976 6316
rect 16028 6332 16080 6384
rect 16672 6307 16724 6316
rect 15476 6196 15528 6248
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 17316 6264 17368 6316
rect 17960 6264 18012 6316
rect 19800 6400 19852 6452
rect 18236 6332 18288 6384
rect 18512 6307 18564 6316
rect 16580 6196 16632 6248
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 19524 6307 19576 6316
rect 19524 6273 19533 6307
rect 19533 6273 19567 6307
rect 19567 6273 19576 6307
rect 19524 6264 19576 6273
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 18696 6196 18748 6248
rect 11980 6128 12032 6180
rect 14188 6128 14240 6180
rect 14464 6128 14516 6180
rect 14924 6128 14976 6180
rect 20168 6128 20220 6180
rect 12348 6060 12400 6112
rect 13728 6060 13780 6112
rect 14004 6060 14056 6112
rect 15016 6060 15068 6112
rect 15200 6060 15252 6112
rect 16304 6060 16356 6112
rect 16396 6060 16448 6112
rect 17132 6060 17184 6112
rect 18420 6060 18472 6112
rect 20076 6060 20128 6112
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 4338 5958 4390 6010
rect 4402 5958 4454 6010
rect 4466 5958 4518 6010
rect 4530 5958 4582 6010
rect 4594 5958 4646 6010
rect 11116 5958 11168 6010
rect 11180 5958 11232 6010
rect 11244 5958 11296 6010
rect 11308 5958 11360 6010
rect 11372 5958 11424 6010
rect 17893 5958 17945 6010
rect 17957 5958 18009 6010
rect 18021 5958 18073 6010
rect 18085 5958 18137 6010
rect 18149 5958 18201 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 4988 5899 5040 5908
rect 4988 5865 4997 5899
rect 4997 5865 5031 5899
rect 5031 5865 5040 5899
rect 4988 5856 5040 5865
rect 5264 5856 5316 5908
rect 7472 5856 7524 5908
rect 9312 5856 9364 5908
rect 16764 5856 16816 5908
rect 17224 5856 17276 5908
rect 18420 5899 18472 5908
rect 2504 5788 2556 5840
rect 2964 5720 3016 5772
rect 5172 5788 5224 5840
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 3792 5652 3844 5704
rect 5264 5720 5316 5772
rect 5356 5720 5408 5772
rect 9588 5788 9640 5840
rect 9680 5788 9732 5840
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 18696 5899 18748 5908
rect 18696 5865 18705 5899
rect 18705 5865 18739 5899
rect 18739 5865 18748 5899
rect 18696 5856 18748 5865
rect 19248 5856 19300 5908
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 4804 5695 4856 5704
rect 4804 5661 4818 5695
rect 4818 5661 4852 5695
rect 4852 5661 4856 5695
rect 6276 5695 6328 5704
rect 4804 5652 4856 5661
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 7472 5652 7524 5704
rect 7656 5652 7708 5704
rect 8576 5720 8628 5772
rect 9312 5720 9364 5772
rect 9956 5720 10008 5772
rect 10600 5720 10652 5772
rect 12716 5763 12768 5772
rect 3700 5584 3752 5636
rect 3240 5516 3292 5568
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 4896 5584 4948 5636
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 5356 5516 5408 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 7656 5516 7708 5568
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 9496 5584 9548 5636
rect 10416 5652 10468 5704
rect 10968 5652 11020 5704
rect 11060 5652 11112 5704
rect 11704 5652 11756 5704
rect 11980 5652 12032 5704
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 13820 5720 13872 5772
rect 14372 5720 14424 5772
rect 15016 5720 15068 5772
rect 13268 5652 13320 5704
rect 14096 5652 14148 5704
rect 14464 5695 14516 5704
rect 10692 5584 10744 5636
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 16028 5652 16080 5704
rect 16304 5695 16356 5704
rect 16304 5661 16313 5695
rect 16313 5661 16347 5695
rect 16347 5661 16356 5695
rect 16304 5652 16356 5661
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 17592 5695 17644 5704
rect 16580 5652 16632 5661
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 20628 5788 20680 5840
rect 18604 5720 18656 5772
rect 20260 5720 20312 5772
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 20352 5652 20404 5704
rect 9956 5516 10008 5568
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 18696 5584 18748 5636
rect 12164 5516 12216 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 13636 5516 13688 5568
rect 17040 5516 17092 5568
rect 18880 5516 18932 5568
rect 20168 5516 20220 5568
rect 7727 5414 7779 5466
rect 7791 5414 7843 5466
rect 7855 5414 7907 5466
rect 7919 5414 7971 5466
rect 7983 5414 8035 5466
rect 14504 5414 14556 5466
rect 14568 5414 14620 5466
rect 14632 5414 14684 5466
rect 14696 5414 14748 5466
rect 14760 5414 14812 5466
rect 3700 5312 3752 5364
rect 6368 5312 6420 5364
rect 9036 5312 9088 5364
rect 9220 5312 9272 5364
rect 1584 5244 1636 5296
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4160 5176 4212 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 7380 5244 7432 5296
rect 5356 5176 5408 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 7748 5176 7800 5228
rect 6920 5108 6972 5160
rect 9680 5244 9732 5296
rect 9864 5287 9916 5296
rect 9864 5253 9873 5287
rect 9873 5253 9907 5287
rect 9907 5253 9916 5287
rect 9864 5244 9916 5253
rect 9128 5176 9180 5228
rect 9220 5176 9272 5228
rect 7656 5083 7708 5092
rect 7656 5049 7665 5083
rect 7665 5049 7699 5083
rect 7699 5049 7708 5083
rect 7656 5040 7708 5049
rect 7840 5040 7892 5092
rect 9864 5108 9916 5160
rect 9956 5108 10008 5160
rect 10600 5108 10652 5160
rect 9588 5040 9640 5092
rect 11060 5312 11112 5364
rect 12624 5312 12676 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 13728 5355 13780 5364
rect 13728 5321 13737 5355
rect 13737 5321 13771 5355
rect 13771 5321 13780 5355
rect 13728 5312 13780 5321
rect 11612 5244 11664 5296
rect 11520 5176 11572 5228
rect 12072 5244 12124 5296
rect 14372 5244 14424 5296
rect 12532 5176 12584 5228
rect 13912 5176 13964 5228
rect 13452 5108 13504 5160
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 14924 5176 14976 5228
rect 16212 5244 16264 5296
rect 17040 5355 17092 5364
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 18696 5312 18748 5364
rect 20352 5355 20404 5364
rect 17684 5176 17736 5228
rect 19064 5244 19116 5296
rect 12348 5040 12400 5092
rect 14188 5040 14240 5092
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 7012 4972 7064 5024
rect 7288 4972 7340 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 9680 4972 9732 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13636 4972 13688 5024
rect 16212 5108 16264 5160
rect 17500 5108 17552 5160
rect 18328 5108 18380 5160
rect 20352 5321 20361 5355
rect 20361 5321 20395 5355
rect 20395 5321 20404 5355
rect 20352 5312 20404 5321
rect 19432 5244 19484 5296
rect 19156 5108 19208 5160
rect 17592 5040 17644 5092
rect 18512 5040 18564 5092
rect 14372 4972 14424 5024
rect 15200 4972 15252 5024
rect 4338 4870 4390 4922
rect 4402 4870 4454 4922
rect 4466 4870 4518 4922
rect 4530 4870 4582 4922
rect 4594 4870 4646 4922
rect 11116 4870 11168 4922
rect 11180 4870 11232 4922
rect 11244 4870 11296 4922
rect 11308 4870 11360 4922
rect 11372 4870 11424 4922
rect 17893 4870 17945 4922
rect 17957 4870 18009 4922
rect 18021 4870 18073 4922
rect 18085 4870 18137 4922
rect 18149 4870 18201 4922
rect 4896 4768 4948 4820
rect 6368 4768 6420 4820
rect 9404 4768 9456 4820
rect 9588 4768 9640 4820
rect 16212 4768 16264 4820
rect 17224 4768 17276 4820
rect 18512 4768 18564 4820
rect 19800 4768 19852 4820
rect 5816 4700 5868 4752
rect 9036 4700 9088 4752
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1768 4564 1820 4616
rect 2688 4564 2740 4616
rect 3700 4564 3752 4616
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 2596 4428 2648 4480
rect 3884 4428 3936 4480
rect 4712 4564 4764 4616
rect 5356 4564 5408 4616
rect 5632 4564 5684 4616
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6828 4564 6880 4616
rect 7748 4564 7800 4616
rect 7012 4496 7064 4548
rect 7840 4496 7892 4548
rect 8208 4539 8260 4548
rect 8208 4505 8217 4539
rect 8217 4505 8251 4539
rect 8251 4505 8260 4539
rect 8208 4496 8260 4505
rect 8852 4496 8904 4548
rect 9588 4564 9640 4616
rect 10048 4632 10100 4684
rect 10508 4700 10560 4752
rect 12624 4632 12676 4684
rect 5080 4428 5132 4480
rect 6920 4428 6972 4480
rect 7104 4428 7156 4480
rect 9588 4428 9640 4480
rect 9772 4496 9824 4548
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 11704 4564 11756 4616
rect 10692 4496 10744 4548
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12256 4607 12308 4616
rect 12072 4564 12124 4573
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 12992 4564 13044 4616
rect 13360 4564 13412 4616
rect 12808 4496 12860 4548
rect 15200 4564 15252 4616
rect 17684 4700 17736 4752
rect 16488 4632 16540 4684
rect 17408 4632 17460 4684
rect 18604 4632 18656 4684
rect 16672 4564 16724 4616
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 16580 4496 16632 4548
rect 17868 4564 17920 4616
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19340 4607 19392 4616
rect 19340 4573 19350 4607
rect 19350 4573 19384 4607
rect 19384 4573 19392 4607
rect 19340 4564 19392 4573
rect 19432 4496 19484 4548
rect 19616 4539 19668 4548
rect 19616 4505 19625 4539
rect 19625 4505 19659 4539
rect 19659 4505 19668 4539
rect 19616 4496 19668 4505
rect 13820 4428 13872 4480
rect 15200 4428 15252 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 19156 4428 19208 4480
rect 20720 4539 20772 4548
rect 20720 4505 20729 4539
rect 20729 4505 20763 4539
rect 20763 4505 20772 4539
rect 20720 4496 20772 4505
rect 7727 4326 7779 4378
rect 7791 4326 7843 4378
rect 7855 4326 7907 4378
rect 7919 4326 7971 4378
rect 7983 4326 8035 4378
rect 14504 4326 14556 4378
rect 14568 4326 14620 4378
rect 14632 4326 14684 4378
rect 14696 4326 14748 4378
rect 14760 4326 14812 4378
rect 5540 4224 5592 4276
rect 7288 4224 7340 4276
rect 9036 4224 9088 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 10876 4224 10928 4276
rect 15936 4267 15988 4276
rect 2596 4199 2648 4208
rect 2596 4165 2605 4199
rect 2605 4165 2639 4199
rect 2639 4165 2648 4199
rect 2596 4156 2648 4165
rect 3700 4156 3752 4208
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 5908 4156 5960 4208
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4988 4131 5040 4140
rect 2872 4020 2924 4072
rect 4252 4020 4304 4072
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 6184 4088 6236 4140
rect 6736 4156 6788 4208
rect 8300 4156 8352 4208
rect 10784 4199 10836 4208
rect 10784 4165 10793 4199
rect 10793 4165 10827 4199
rect 10827 4165 10836 4199
rect 10784 4156 10836 4165
rect 12900 4199 12952 4208
rect 5080 4020 5132 4072
rect 3976 3952 4028 4004
rect 4712 3952 4764 4004
rect 5448 3952 5500 4004
rect 8024 4088 8076 4140
rect 10048 4131 10100 4140
rect 9772 4020 9824 4072
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 10324 4088 10376 4140
rect 12900 4165 12909 4199
rect 12909 4165 12943 4199
rect 12943 4165 12952 4199
rect 12900 4156 12952 4165
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 16580 4224 16632 4276
rect 12624 4131 12676 4140
rect 11704 4020 11756 4072
rect 12072 4020 12124 4072
rect 7288 3952 7340 4004
rect 9404 3952 9456 4004
rect 2780 3884 2832 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 4068 3884 4120 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6644 3884 6696 3936
rect 8300 3884 8352 3936
rect 9036 3884 9088 3936
rect 9128 3884 9180 3936
rect 10692 3884 10744 3936
rect 11520 3952 11572 4004
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 13268 4088 13320 4140
rect 13452 4088 13504 4140
rect 15108 4088 15160 4140
rect 15844 4088 15896 4140
rect 15936 4088 15988 4140
rect 16856 4156 16908 4208
rect 17408 4224 17460 4276
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17868 4156 17920 4208
rect 19156 4224 19208 4276
rect 14740 4020 14792 4072
rect 16580 4020 16632 4072
rect 11612 3884 11664 3936
rect 11796 3884 11848 3936
rect 19616 4156 19668 4208
rect 18236 4088 18288 4140
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 19708 4088 19760 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 19340 4020 19392 4072
rect 20812 3952 20864 4004
rect 12992 3884 13044 3936
rect 13084 3884 13136 3936
rect 15200 3884 15252 3936
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 20076 3884 20128 3936
rect 21364 3884 21416 3936
rect 4338 3782 4390 3834
rect 4402 3782 4454 3834
rect 4466 3782 4518 3834
rect 4530 3782 4582 3834
rect 4594 3782 4646 3834
rect 11116 3782 11168 3834
rect 11180 3782 11232 3834
rect 11244 3782 11296 3834
rect 11308 3782 11360 3834
rect 11372 3782 11424 3834
rect 17893 3782 17945 3834
rect 17957 3782 18009 3834
rect 18021 3782 18073 3834
rect 18085 3782 18137 3834
rect 18149 3782 18201 3834
rect 2964 3680 3016 3732
rect 3700 3680 3752 3732
rect 5540 3680 5592 3732
rect 6460 3680 6512 3732
rect 7656 3680 7708 3732
rect 9772 3680 9824 3732
rect 10140 3680 10192 3732
rect 10416 3723 10468 3732
rect 10416 3689 10425 3723
rect 10425 3689 10459 3723
rect 10459 3689 10468 3723
rect 10416 3680 10468 3689
rect 11704 3723 11756 3732
rect 11704 3689 11713 3723
rect 11713 3689 11747 3723
rect 11747 3689 11756 3723
rect 11704 3680 11756 3689
rect 12164 3680 12216 3732
rect 12624 3680 12676 3732
rect 14280 3680 14332 3732
rect 15292 3680 15344 3732
rect 16580 3680 16632 3732
rect 17776 3680 17828 3732
rect 18420 3723 18472 3732
rect 18420 3689 18429 3723
rect 18429 3689 18463 3723
rect 18463 3689 18472 3723
rect 18420 3680 18472 3689
rect 3976 3476 4028 3528
rect 4252 3612 4304 3664
rect 4344 3612 4396 3664
rect 5356 3612 5408 3664
rect 5172 3544 5224 3596
rect 4528 3476 4580 3528
rect 5724 3544 5776 3596
rect 1492 3408 1544 3460
rect 3056 3451 3108 3460
rect 3056 3417 3065 3451
rect 3065 3417 3099 3451
rect 3099 3417 3108 3451
rect 3056 3408 3108 3417
rect 4160 3451 4212 3460
rect 4160 3417 4169 3451
rect 4169 3417 4203 3451
rect 4203 3417 4212 3451
rect 4160 3408 4212 3417
rect 4344 3408 4396 3460
rect 5632 3476 5684 3528
rect 6184 3476 6236 3528
rect 6368 3476 6420 3528
rect 6920 3612 6972 3664
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7288 3519 7340 3528
rect 7012 3476 7064 3485
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7380 3476 7432 3528
rect 8024 3476 8076 3528
rect 9680 3544 9732 3596
rect 10048 3544 10100 3596
rect 9312 3476 9364 3528
rect 10232 3476 10284 3528
rect 10508 3476 10560 3528
rect 12072 3544 12124 3596
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 12348 3544 12400 3553
rect 13268 3612 13320 3664
rect 13912 3612 13964 3664
rect 15016 3612 15068 3664
rect 16672 3612 16724 3664
rect 18604 3612 18656 3664
rect 17224 3544 17276 3596
rect 17868 3544 17920 3596
rect 19340 3544 19392 3596
rect 20 3340 72 3392
rect 2228 3340 2280 3392
rect 3976 3340 4028 3392
rect 10876 3451 10928 3460
rect 10876 3417 10911 3451
rect 10911 3417 10928 3451
rect 10876 3408 10928 3417
rect 4528 3340 4580 3392
rect 4804 3340 4856 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 7012 3340 7064 3392
rect 9680 3340 9732 3392
rect 10140 3340 10192 3392
rect 11980 3476 12032 3528
rect 12900 3476 12952 3528
rect 13636 3476 13688 3528
rect 14832 3476 14884 3528
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 15936 3476 15988 3528
rect 11612 3408 11664 3460
rect 17960 3476 18012 3528
rect 18144 3476 18196 3528
rect 19708 3476 19760 3528
rect 16396 3451 16448 3460
rect 16396 3417 16405 3451
rect 16405 3417 16439 3451
rect 16439 3417 16448 3451
rect 16396 3408 16448 3417
rect 19524 3451 19576 3460
rect 19524 3417 19533 3451
rect 19533 3417 19567 3451
rect 19567 3417 19576 3451
rect 19524 3408 19576 3417
rect 19984 3451 20036 3460
rect 19984 3417 19993 3451
rect 19993 3417 20027 3451
rect 20027 3417 20036 3451
rect 19984 3408 20036 3417
rect 21916 3408 21968 3460
rect 12164 3340 12216 3392
rect 13268 3340 13320 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 15660 3340 15712 3392
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 17500 3340 17552 3392
rect 17868 3340 17920 3392
rect 18328 3340 18380 3392
rect 7727 3238 7779 3290
rect 7791 3238 7843 3290
rect 7855 3238 7907 3290
rect 7919 3238 7971 3290
rect 7983 3238 8035 3290
rect 14504 3238 14556 3290
rect 14568 3238 14620 3290
rect 14632 3238 14684 3290
rect 14696 3238 14748 3290
rect 14760 3238 14812 3290
rect 1492 3179 1544 3188
rect 1492 3145 1501 3179
rect 1501 3145 1535 3179
rect 1535 3145 1544 3179
rect 1492 3136 1544 3145
rect 2136 3068 2188 3120
rect 3148 3068 3200 3120
rect 3792 3068 3844 3120
rect 2688 3000 2740 3052
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 5356 3136 5408 3188
rect 6184 3136 6236 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 8392 3136 8444 3188
rect 9588 3179 9640 3188
rect 7288 3068 7340 3120
rect 5540 3000 5592 3052
rect 5632 3000 5684 3052
rect 572 2864 624 2916
rect 1124 2796 1176 2848
rect 3516 2864 3568 2916
rect 4896 2932 4948 2984
rect 4988 2932 5040 2984
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 8300 3000 8352 3052
rect 8208 2864 8260 2916
rect 3056 2796 3108 2848
rect 8576 2932 8628 2984
rect 9588 3145 9597 3179
rect 9597 3145 9631 3179
rect 9631 3145 9640 3179
rect 9588 3136 9640 3145
rect 10508 3179 10560 3188
rect 10508 3145 10517 3179
rect 10517 3145 10551 3179
rect 10551 3145 10560 3179
rect 10508 3136 10560 3145
rect 12256 3136 12308 3188
rect 12440 3136 12492 3188
rect 12532 3136 12584 3188
rect 14096 3136 14148 3188
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 18236 3136 18288 3188
rect 9772 3068 9824 3120
rect 10048 3068 10100 3120
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 10876 3068 10928 3120
rect 11980 3068 12032 3120
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9680 3000 9732 3052
rect 12808 3068 12860 3120
rect 14372 3068 14424 3120
rect 12716 3043 12768 3052
rect 9864 2932 9916 2984
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 13360 3043 13412 3052
rect 13360 3009 13369 3043
rect 13369 3009 13403 3043
rect 13403 3009 13412 3043
rect 13360 3000 13412 3009
rect 13636 3000 13688 3052
rect 17408 3068 17460 3120
rect 15016 3000 15068 3052
rect 8760 2864 8812 2916
rect 12164 2864 12216 2916
rect 16120 2932 16172 2984
rect 16304 2932 16356 2984
rect 17132 3000 17184 3052
rect 16856 2932 16908 2984
rect 18236 3000 18288 3052
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 20260 3000 20312 3052
rect 18420 2932 18472 2984
rect 12440 2864 12492 2916
rect 16396 2796 16448 2848
rect 4338 2694 4390 2746
rect 4402 2694 4454 2746
rect 4466 2694 4518 2746
rect 4530 2694 4582 2746
rect 4594 2694 4646 2746
rect 11116 2694 11168 2746
rect 11180 2694 11232 2746
rect 11244 2694 11296 2746
rect 11308 2694 11360 2746
rect 11372 2694 11424 2746
rect 17893 2694 17945 2746
rect 17957 2694 18009 2746
rect 18021 2694 18073 2746
rect 18085 2694 18137 2746
rect 18149 2694 18201 2746
rect 4160 2524 4212 2576
rect 8484 2524 8536 2576
rect 9312 2592 9364 2644
rect 12256 2592 12308 2644
rect 14188 2592 14240 2644
rect 11612 2524 11664 2576
rect 8944 2456 8996 2508
rect 12072 2456 12124 2508
rect 13360 2456 13412 2508
rect 1676 2388 1728 2440
rect 5356 2388 5408 2440
rect 6460 2388 6512 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 11796 2388 11848 2440
rect 16764 2592 16816 2644
rect 17684 2592 17736 2644
rect 19156 2592 19208 2644
rect 15568 2524 15620 2576
rect 16948 2456 17000 2508
rect 17132 2456 17184 2508
rect 18604 2456 18656 2508
rect 16580 2388 16632 2440
rect 18972 2388 19024 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 2412 2320 2464 2372
rect 2964 2320 3016 2372
rect 5908 2320 5960 2372
rect 4344 2295 4396 2304
rect 4344 2261 4353 2295
rect 4353 2261 4387 2295
rect 4387 2261 4396 2295
rect 4344 2252 4396 2261
rect 8300 2320 8352 2372
rect 12532 2320 12584 2372
rect 15476 2320 15528 2372
rect 17316 2320 17368 2372
rect 13176 2252 13228 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 18788 2252 18840 2304
rect 7727 2150 7779 2202
rect 7791 2150 7843 2202
rect 7855 2150 7907 2202
rect 7919 2150 7971 2202
rect 7983 2150 8035 2202
rect 14504 2150 14556 2202
rect 14568 2150 14620 2202
rect 14632 2150 14684 2202
rect 14696 2150 14748 2202
rect 14760 2150 14812 2202
rect 4344 2048 4396 2100
rect 19064 2048 19116 2100
rect 7564 1980 7616 2032
rect 13360 1980 13412 2032
rect 16764 1980 16816 2032
rect 19892 1980 19944 2032
<< metal2 >>
rect 570 23911 626 24711
rect 1122 23911 1178 24711
rect 1674 23911 1730 24711
rect 2226 23911 2282 24711
rect 2778 23911 2834 24711
rect 3146 24576 3202 24585
rect 3146 24511 3202 24520
rect 584 21146 612 23911
rect 572 21140 624 21146
rect 572 21082 624 21088
rect 1136 20942 1164 23911
rect 1124 20936 1176 20942
rect 1124 20878 1176 20884
rect 1582 20224 1638 20233
rect 1582 20159 1638 20168
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19417 1440 19790
rect 1596 19514 1624 20159
rect 1688 19990 1716 23911
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1872 21622 1900 22063
rect 1860 21616 1912 21622
rect 1860 21558 1912 21564
rect 1768 21412 1820 21418
rect 1768 21354 1820 21360
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1398 19408 1454 19417
rect 1688 19378 1716 19790
rect 1398 19343 1454 19352
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1216 19304 1268 19310
rect 1216 19246 1268 19252
rect 1228 10169 1256 19246
rect 1308 16584 1360 16590
rect 1308 16526 1360 16532
rect 1320 12220 1348 16526
rect 1504 16250 1532 19314
rect 1674 18592 1730 18601
rect 1674 18527 1730 18536
rect 1688 18426 1716 18527
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17338 1624 18226
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1780 15638 1808 21354
rect 2240 21078 2268 23911
rect 2792 23882 2820 23911
rect 2700 23854 2820 23882
rect 2318 22944 2374 22953
rect 2318 22879 2374 22888
rect 2228 21072 2280 21078
rect 2228 21014 2280 21020
rect 2332 20602 2360 22879
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2148 18766 2176 19314
rect 2240 18970 2268 20402
rect 2318 19408 2374 19417
rect 2318 19343 2320 19352
rect 2372 19343 2374 19352
rect 2320 19314 2372 19320
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1872 17513 1900 17546
rect 1952 17536 2004 17542
rect 1858 17504 1914 17513
rect 1952 17478 2004 17484
rect 1858 17439 1914 17448
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 13977 1716 14282
rect 1674 13968 1730 13977
rect 1492 13932 1544 13938
rect 1674 13903 1730 13912
rect 1492 13874 1544 13880
rect 1504 12442 1532 13874
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13161 1624 13670
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1400 12232 1452 12238
rect 1320 12192 1400 12220
rect 1400 12174 1452 12180
rect 1214 10160 1270 10169
rect 1214 10095 1270 10104
rect 1412 9586 1440 12174
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1504 9450 1532 11698
rect 1584 11552 1636 11558
rect 1582 11520 1584 11529
rect 1636 11520 1638 11529
rect 1582 11455 1638 11464
rect 1584 10464 1636 10470
rect 1582 10432 1584 10441
rect 1636 10432 1638 10441
rect 1582 10367 1638 10376
rect 1780 10010 1808 14350
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 12345 1900 12786
rect 1858 12336 1914 12345
rect 1858 12271 1914 12280
rect 1964 10690 1992 17478
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16590 2084 17138
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2240 16046 2268 18770
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2424 17746 2452 18294
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2516 17338 2544 20810
rect 2700 20398 2728 23854
rect 2778 23760 2834 23769
rect 2778 23695 2834 23704
rect 2792 22030 2820 23695
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 3160 21554 3188 24511
rect 3514 23911 3570 24711
rect 4066 23911 4122 24711
rect 4618 23911 4674 24711
rect 5170 23911 5226 24711
rect 5906 23911 5962 24711
rect 6458 23911 6514 24711
rect 7010 23911 7066 24711
rect 7562 23911 7618 24711
rect 8298 23911 8354 24711
rect 8850 23911 8906 24711
rect 9402 23911 9458 24711
rect 9954 23911 10010 24711
rect 10690 23911 10746 24711
rect 10796 23990 11008 24018
rect 3528 22030 3556 23911
rect 4080 22098 4108 23911
rect 4632 22522 4660 23911
rect 4632 22494 4752 22522
rect 4338 22332 4646 22352
rect 4338 22330 4344 22332
rect 4400 22330 4424 22332
rect 4480 22330 4504 22332
rect 4560 22330 4584 22332
rect 4640 22330 4646 22332
rect 4400 22278 4402 22330
rect 4582 22278 4584 22330
rect 4338 22276 4344 22278
rect 4400 22276 4424 22278
rect 4480 22276 4504 22278
rect 4560 22276 4584 22278
rect 4640 22276 4646 22278
rect 4338 22256 4646 22276
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3068 20534 3096 21286
rect 3238 21040 3294 21049
rect 3238 20975 3294 20984
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 19786 2912 20266
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2884 19310 2912 19722
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2976 18970 3004 20198
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 3068 19310 3096 19722
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19514 3188 19654
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2608 18426 2636 18702
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2976 17678 3004 18906
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 3252 16590 3280 20975
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 18426 3464 18566
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3344 17678 3372 18158
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 17241 3372 17614
rect 3330 17232 3386 17241
rect 3330 17167 3386 17176
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2228 16040 2280 16046
rect 2700 16017 2728 16390
rect 2228 15982 2280 15988
rect 2686 16008 2742 16017
rect 2056 15706 2084 15982
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2148 13394 2176 13670
rect 2240 13394 2268 15982
rect 2686 15943 2742 15952
rect 2792 15881 2820 16526
rect 3332 16108 3384 16114
rect 3252 16068 3332 16096
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2424 13938 2452 14486
rect 2516 14414 2544 15370
rect 2608 15026 2636 15506
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2608 14822 2636 14962
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14414 2636 14758
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2608 14226 2636 14350
rect 2516 14198 2636 14226
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 10810 2084 12174
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 1964 10662 2084 10690
rect 2148 10674 2176 11834
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10742 2268 11018
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 1676 9988 1728 9994
rect 1780 9982 1900 10010
rect 1676 9930 1728 9936
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1688 8401 1716 9930
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 9625 1808 9862
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 1872 9518 1900 9982
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1674 7984 1730 7993
rect 1674 7919 1730 7928
rect 1688 7886 1716 7919
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 6656 1636 6662
rect 1780 6633 1808 9454
rect 1952 8832 2004 8838
rect 1950 8800 1952 8809
rect 2004 8800 2006 8809
rect 1950 8735 2006 8744
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7818 1992 8230
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 6905 1900 7346
rect 2056 6914 2084 10662
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2332 9874 2360 13126
rect 2516 11150 2544 14198
rect 2700 13190 2728 15438
rect 2792 15065 2820 15438
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2884 14958 2912 15982
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2976 15162 3004 15438
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14414 2912 14894
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2792 12918 2820 13738
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2884 12850 2912 13466
rect 2976 12850 3004 13942
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2424 10062 2452 11086
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2516 10266 2544 10746
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10062 2636 12038
rect 2700 11898 2728 12582
rect 3068 12306 3096 15846
rect 3252 15366 3280 16068
rect 3332 16050 3384 16056
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15094 3280 15302
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3514 15056 3570 15065
rect 3252 14618 3280 15030
rect 3514 14991 3570 15000
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3160 13530 3188 13874
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3252 12850 3280 13738
rect 3344 13326 3372 14010
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3436 13530 3464 13874
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 12442 3188 12718
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 12306 3280 12786
rect 3436 12782 3464 13262
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3528 12628 3556 14991
rect 3436 12600 3556 12628
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2700 11762 2728 11834
rect 2884 11762 2912 12038
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11642 2912 11698
rect 2700 11614 2912 11642
rect 2700 11354 2728 11614
rect 2872 11552 2924 11558
rect 2976 11540 3004 12106
rect 2924 11512 3004 11540
rect 2872 11494 2924 11500
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2700 11150 2728 11290
rect 2884 11218 2912 11494
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2332 9846 2452 9874
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2148 8634 2176 9318
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2148 7954 2176 8570
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2056 6905 2268 6914
rect 1858 6896 1914 6905
rect 2056 6896 2282 6905
rect 2056 6886 2226 6896
rect 1858 6831 1914 6840
rect 2226 6831 2282 6840
rect 2332 6798 2360 7686
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2044 6656 2096 6662
rect 1584 6598 1636 6604
rect 1766 6624 1822 6633
rect 1596 5302 1624 6598
rect 2044 6598 2096 6604
rect 1766 6559 1822 6568
rect 1780 6322 1808 6559
rect 2056 6458 2084 6598
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2332 6322 2360 6734
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1780 4622 1808 6258
rect 2136 6112 2188 6118
rect 1950 6080 2006 6089
rect 2136 6054 2188 6060
rect 1950 6015 2006 6024
rect 1964 5914 1992 6015
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1860 5704 1912 5710
rect 1858 5672 1860 5681
rect 1912 5672 1914 5681
rect 1858 5607 1914 5616
rect 2042 5264 2098 5273
rect 2042 5199 2044 5208
rect 2096 5199 2098 5208
rect 2044 5170 2096 5176
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1412 4457 1440 4558
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 20 3392 72 3398
rect 20 3334 72 3340
rect 32 800 60 3334
rect 1504 3194 1532 3402
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 2148 3126 2176 6054
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 584 800 612 2858
rect 1124 2848 1176 2854
rect 1124 2790 1176 2796
rect 1136 800 1164 2790
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 800 1716 2382
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 921 1900 2314
rect 1858 912 1914 921
rect 1858 847 1914 856
rect 2240 800 2268 3334
rect 2424 2378 2452 9846
rect 2700 9586 2728 10950
rect 2792 10742 2820 11086
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2884 10062 2912 11154
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 10674 3372 11018
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2976 9654 3004 10406
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2700 8974 2728 9522
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2516 8430 2544 8570
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2516 7886 2544 8366
rect 2792 7954 2820 8434
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2884 7886 2912 8502
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2516 6390 2544 7822
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2516 5846 2544 6326
rect 2608 6322 2636 6598
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2884 6254 2912 6938
rect 2976 6322 3004 9590
rect 3436 9586 3464 12600
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2976 5914 3004 6122
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2608 4214 2636 4422
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2700 3058 2728 4558
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2792 2553 2820 3878
rect 2778 2544 2834 2553
rect 2778 2479 2834 2488
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2884 1737 2912 4014
rect 2976 3738 3004 5714
rect 3068 5234 3096 9522
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3620 8922 3648 21898
rect 4338 21244 4646 21264
rect 4338 21242 4344 21244
rect 4400 21242 4424 21244
rect 4480 21242 4504 21244
rect 4560 21242 4584 21244
rect 4640 21242 4646 21244
rect 4400 21190 4402 21242
rect 4582 21190 4584 21242
rect 4338 21188 4344 21190
rect 4400 21188 4424 21190
rect 4480 21188 4504 21190
rect 4560 21188 4584 21190
rect 4640 21188 4646 21190
rect 4338 21168 4646 21188
rect 4724 21146 4752 22494
rect 4896 21616 4948 21622
rect 4896 21558 4948 21564
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4172 20602 4200 20742
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4264 20534 4292 20742
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3896 19446 3924 20402
rect 3976 20256 4028 20262
rect 4356 20244 4384 20946
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 3976 20198 4028 20204
rect 4264 20216 4384 20244
rect 4712 20256 4764 20262
rect 3884 19440 3936 19446
rect 3712 19400 3884 19428
rect 3712 17202 3740 19400
rect 3884 19382 3936 19388
rect 3988 19394 4016 20198
rect 4264 19938 4292 20216
rect 4712 20198 4764 20204
rect 4338 20156 4646 20176
rect 4338 20154 4344 20156
rect 4400 20154 4424 20156
rect 4480 20154 4504 20156
rect 4560 20154 4584 20156
rect 4640 20154 4646 20156
rect 4400 20102 4402 20154
rect 4582 20102 4584 20154
rect 4338 20100 4344 20102
rect 4400 20100 4424 20102
rect 4480 20100 4504 20102
rect 4560 20100 4584 20102
rect 4640 20100 4646 20102
rect 4338 20080 4646 20100
rect 4724 20058 4752 20198
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4264 19922 4384 19938
rect 4264 19916 4396 19922
rect 4264 19910 4344 19916
rect 4344 19858 4396 19864
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4080 19514 4108 19654
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3988 19366 4108 19394
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3882 19272 3938 19281
rect 3804 18766 3832 19246
rect 3882 19207 3884 19216
rect 3936 19207 3938 19216
rect 3884 19178 3936 19184
rect 4080 19174 4108 19366
rect 4160 19304 4212 19310
rect 4264 19281 4292 19654
rect 4160 19246 4212 19252
rect 4250 19272 4306 19281
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 3804 16250 3832 18702
rect 3896 17542 3924 18702
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3988 17746 4016 18226
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3896 16522 3924 17478
rect 3988 16572 4016 17682
rect 4080 17649 4108 19110
rect 4172 18970 4200 19246
rect 4250 19207 4306 19216
rect 4356 19156 4384 19858
rect 4540 19378 4568 19858
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4264 19128 4384 19156
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4264 18170 4292 19128
rect 4338 19068 4646 19088
rect 4338 19066 4344 19068
rect 4400 19066 4424 19068
rect 4480 19066 4504 19068
rect 4560 19066 4584 19068
rect 4640 19066 4646 19068
rect 4400 19014 4402 19066
rect 4582 19014 4584 19066
rect 4338 19012 4344 19014
rect 4400 19012 4424 19014
rect 4480 19012 4504 19014
rect 4560 19012 4584 19014
rect 4640 19012 4646 19014
rect 4338 18992 4646 19012
rect 4172 18142 4292 18170
rect 4172 17746 4200 18142
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4066 17640 4122 17649
rect 4066 17575 4122 17584
rect 4080 17066 4108 17575
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 17338 4200 17478
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4264 17202 4292 18022
rect 4338 17980 4646 18000
rect 4338 17978 4344 17980
rect 4400 17978 4424 17980
rect 4480 17978 4504 17980
rect 4560 17978 4584 17980
rect 4640 17978 4646 17980
rect 4400 17926 4402 17978
rect 4582 17926 4584 17978
rect 4338 17924 4344 17926
rect 4400 17924 4424 17926
rect 4480 17924 4504 17926
rect 4560 17924 4584 17926
rect 4640 17924 4646 17926
rect 4338 17904 4646 17924
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4338 16892 4646 16912
rect 4338 16890 4344 16892
rect 4400 16890 4424 16892
rect 4480 16890 4504 16892
rect 4560 16890 4584 16892
rect 4640 16890 4646 16892
rect 4400 16838 4402 16890
rect 4582 16838 4584 16890
rect 4338 16836 4344 16838
rect 4400 16836 4424 16838
rect 4480 16836 4504 16838
rect 4560 16836 4584 16838
rect 4640 16836 4646 16838
rect 4338 16816 4646 16836
rect 4066 16688 4122 16697
rect 4122 16646 4200 16674
rect 4066 16623 4122 16632
rect 3988 16544 4108 16572
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 4080 16454 4108 16544
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 4172 16114 4200 16646
rect 4724 16590 4752 19790
rect 4816 19417 4844 20402
rect 4802 19408 4858 19417
rect 4802 19343 4858 19352
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 3804 15706 3832 16050
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 12850 3740 13670
rect 3804 13326 3832 15642
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14006 3924 14214
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3804 12434 3832 12854
rect 3712 12406 3832 12434
rect 3712 11286 3740 12406
rect 3792 12368 3844 12374
rect 3988 12345 4016 15574
rect 4172 13870 4200 15914
rect 4264 14618 4292 16526
rect 4816 16402 4844 19343
rect 4908 16454 4936 21558
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 5000 19378 5028 21014
rect 5080 20868 5132 20874
rect 5080 20810 5132 20816
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5092 18442 5120 20810
rect 5184 19718 5212 23911
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5368 21690 5396 22102
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5368 21486 5396 21626
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5368 20505 5396 20538
rect 5354 20496 5410 20505
rect 5354 20431 5410 20440
rect 5356 20392 5408 20398
rect 5354 20360 5356 20369
rect 5408 20360 5410 20369
rect 5460 20330 5488 21490
rect 5552 20942 5580 21830
rect 5736 20942 5764 22034
rect 5920 22030 5948 23911
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5354 20295 5410 20304
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5460 19854 5488 20266
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5552 19242 5580 20742
rect 5644 19854 5672 20742
rect 5736 20448 5764 20878
rect 5828 20641 5856 20946
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5814 20632 5870 20641
rect 5920 20602 5948 20878
rect 5814 20567 5870 20576
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5816 20460 5868 20466
rect 5736 20420 5816 20448
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5644 19334 5672 19654
rect 5736 19514 5764 20420
rect 5816 20402 5868 20408
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5644 19306 5764 19334
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5000 18414 5120 18442
rect 5000 16794 5028 18414
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 5092 17542 5120 18226
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17338 5120 17478
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5184 17134 5212 18906
rect 5736 18714 5764 19306
rect 5828 18834 5856 19654
rect 5920 19446 5948 19926
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5908 18760 5960 18766
rect 5736 18698 5856 18714
rect 5908 18702 5960 18708
rect 5448 18692 5500 18698
rect 5736 18692 5868 18698
rect 5736 18686 5816 18692
rect 5448 18634 5500 18640
rect 5816 18634 5868 18640
rect 5460 18578 5488 18634
rect 5632 18624 5684 18630
rect 5460 18550 5580 18578
rect 5632 18566 5684 18572
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5184 16794 5212 17070
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 4724 16374 4844 16402
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4338 15804 4646 15824
rect 4338 15802 4344 15804
rect 4400 15802 4424 15804
rect 4480 15802 4504 15804
rect 4560 15802 4584 15804
rect 4640 15802 4646 15804
rect 4400 15750 4402 15802
rect 4582 15750 4584 15802
rect 4338 15748 4344 15750
rect 4400 15748 4424 15750
rect 4480 15748 4504 15750
rect 4560 15748 4584 15750
rect 4640 15748 4646 15750
rect 4338 15728 4646 15748
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 14890 4660 15302
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4338 14716 4646 14736
rect 4338 14714 4344 14716
rect 4400 14714 4424 14716
rect 4480 14714 4504 14716
rect 4560 14714 4584 14716
rect 4640 14714 4646 14716
rect 4400 14662 4402 14714
rect 4582 14662 4584 14714
rect 4338 14660 4344 14662
rect 4400 14660 4424 14662
rect 4480 14660 4504 14662
rect 4560 14660 4584 14662
rect 4640 14660 4646 14662
rect 4338 14640 4646 14660
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4338 13628 4646 13648
rect 4338 13626 4344 13628
rect 4400 13626 4424 13628
rect 4480 13626 4504 13628
rect 4560 13626 4584 13628
rect 4640 13626 4646 13628
rect 4400 13574 4402 13626
rect 4582 13574 4584 13626
rect 4338 13572 4344 13574
rect 4400 13572 4424 13574
rect 4480 13572 4504 13574
rect 4560 13572 4584 13574
rect 4640 13572 4646 13574
rect 4338 13552 4646 13572
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12714 4660 13126
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4338 12540 4646 12560
rect 4338 12538 4344 12540
rect 4400 12538 4424 12540
rect 4480 12538 4504 12540
rect 4560 12538 4584 12540
rect 4640 12538 4646 12540
rect 4400 12486 4402 12538
rect 4582 12486 4584 12538
rect 4338 12484 4344 12486
rect 4400 12484 4424 12486
rect 4480 12484 4504 12486
rect 4560 12484 4584 12486
rect 4640 12484 4646 12486
rect 4338 12464 4646 12484
rect 3792 12310 3844 12316
rect 3974 12336 4030 12345
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3804 10674 3832 12310
rect 3974 12271 4030 12280
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3896 10062 3924 11766
rect 4080 11762 4108 12038
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3988 10810 4016 11698
rect 4080 11150 4108 11698
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4172 10674 4200 11494
rect 4264 11354 4292 11494
rect 4338 11452 4646 11472
rect 4338 11450 4344 11452
rect 4400 11450 4424 11452
rect 4480 11450 4504 11452
rect 4560 11450 4584 11452
rect 4640 11450 4646 11452
rect 4400 11398 4402 11450
rect 4582 11398 4584 11450
rect 4338 11396 4344 11398
rect 4400 11396 4424 11398
rect 4480 11396 4504 11398
rect 4560 11396 4584 11398
rect 4640 11396 4646 11398
rect 4338 11376 4646 11396
rect 4724 11354 4752 16374
rect 4908 16096 4936 16390
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4816 16068 4936 16096
rect 4816 15162 4844 16068
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4816 14822 4844 15098
rect 4908 15094 4936 15914
rect 5000 15570 5028 16186
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 5000 14346 5028 14962
rect 5092 14618 5120 15982
rect 5276 15638 5304 17750
rect 5368 16658 5396 18226
rect 5552 18154 5580 18550
rect 5644 18290 5672 18566
rect 5736 18426 5764 18566
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 18154 5672 18226
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5552 17678 5580 18090
rect 5736 17882 5764 18362
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5920 17762 5948 18702
rect 5644 17734 5948 17762
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5540 17264 5592 17270
rect 5644 17252 5672 17734
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5592 17224 5672 17252
rect 5540 17206 5592 17212
rect 5828 17134 5856 17614
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16114 5764 16390
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5000 13938 5028 14282
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5092 13394 5120 14554
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 13734 5212 14418
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12850 4844 13126
rect 5092 12866 5120 13330
rect 5092 12850 5212 12866
rect 4804 12844 4856 12850
rect 5092 12844 5224 12850
rect 5092 12838 5172 12844
rect 4804 12786 4856 12792
rect 5172 12786 5224 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12306 4936 12582
rect 5276 12306 5304 15574
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14414 5396 14758
rect 5356 14408 5408 14414
rect 5408 14368 5488 14396
rect 5356 14350 5408 14356
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5368 12306 5396 14010
rect 5460 13938 5488 14368
rect 5552 14346 5580 16050
rect 5736 15502 5764 16050
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15162 5764 15302
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5828 15026 5856 15982
rect 6012 15178 6040 21830
rect 6288 21570 6316 21966
rect 6184 21548 6236 21554
rect 6288 21542 6408 21570
rect 6184 21490 6236 21496
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6104 20369 6132 20402
rect 6090 20360 6146 20369
rect 6196 20330 6224 21490
rect 6380 21486 6408 21542
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6380 21128 6408 21422
rect 6288 21100 6408 21128
rect 6288 20806 6316 21100
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6276 20528 6328 20534
rect 6274 20496 6276 20505
rect 6328 20496 6330 20505
rect 6274 20431 6330 20440
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6090 20295 6146 20304
rect 6184 20324 6236 20330
rect 6104 19174 6132 20295
rect 6184 20266 6236 20272
rect 6288 19446 6316 20334
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6380 19334 6408 20810
rect 6472 20058 6500 23911
rect 7024 22094 7052 23911
rect 7024 22066 7144 22094
rect 6644 22024 6696 22030
rect 6564 21984 6644 22012
rect 6564 21554 6592 21984
rect 6644 21966 6696 21972
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6380 19306 6500 19334
rect 6184 19236 6236 19242
rect 6184 19178 6236 19184
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6196 18630 6224 19178
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6380 18290 6408 18770
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6196 17270 6224 17614
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6012 15150 6132 15178
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5724 14816 5776 14822
rect 5722 14784 5724 14793
rect 5776 14784 5778 14793
rect 5722 14719 5778 14728
rect 5828 14618 5856 14962
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5828 14113 5856 14554
rect 5814 14104 5870 14113
rect 5814 14039 5870 14048
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13394 5580 13738
rect 5736 13530 5764 13806
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5460 12850 5488 13194
rect 5828 12918 5856 13194
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5552 12442 5580 12718
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 5276 11676 5304 12242
rect 5368 12186 5396 12242
rect 5368 12158 5488 12186
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11898 5396 12038
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5356 11688 5408 11694
rect 5276 11648 5356 11676
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 10266 4200 10610
rect 4264 10606 4292 11290
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10674 4752 11154
rect 4816 10810 4844 11630
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4338 10364 4646 10384
rect 4338 10362 4344 10364
rect 4400 10362 4424 10364
rect 4480 10362 4504 10364
rect 4560 10362 4584 10364
rect 4640 10362 4646 10364
rect 4400 10310 4402 10362
rect 4582 10310 4584 10362
rect 4338 10308 4344 10310
rect 4400 10308 4424 10310
rect 4480 10308 4504 10310
rect 4560 10308 4584 10310
rect 4640 10308 4646 10310
rect 4338 10288 4646 10308
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 3712 9042 3740 9318
rect 4338 9276 4646 9296
rect 4338 9274 4344 9276
rect 4400 9274 4424 9276
rect 4480 9274 4504 9276
rect 4560 9274 4584 9276
rect 4640 9274 4646 9276
rect 4400 9222 4402 9274
rect 4582 9222 4584 9274
rect 4338 9220 4344 9222
rect 4400 9220 4424 9222
rect 4480 9220 4504 9222
rect 4560 9220 4584 9222
rect 4640 9220 4646 9222
rect 4338 9200 4646 9220
rect 4158 9072 4214 9081
rect 3700 9036 3752 9042
rect 5000 9042 5028 9318
rect 4158 9007 4214 9016
rect 4988 9036 5040 9042
rect 3700 8978 3752 8984
rect 4172 8974 4200 9007
rect 4988 8978 5040 8984
rect 4160 8968 4212 8974
rect 3160 8430 3188 8910
rect 3620 8894 3740 8922
rect 4160 8910 4212 8916
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3514 7984 3570 7993
rect 3514 7919 3570 7928
rect 3528 6866 3556 7919
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 2854 3096 3402
rect 3160 3126 3188 6394
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5234 3280 5510
rect 3620 5234 3648 8774
rect 3712 7857 3740 8894
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3804 8566 3832 8774
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3804 8294 3832 8502
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3896 8090 3924 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7970 4016 8774
rect 4172 8498 4200 8910
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3896 7942 4016 7970
rect 3896 7886 3924 7942
rect 3884 7880 3936 7886
rect 3698 7848 3754 7857
rect 3884 7822 3936 7828
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3698 7783 3754 7792
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3712 7410 3740 7686
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3712 6780 3740 7346
rect 3804 7002 3832 7346
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3792 6792 3844 6798
rect 3712 6752 3792 6780
rect 3792 6734 3844 6740
rect 3804 6322 3832 6734
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5710 3832 6054
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3712 5370 3740 5578
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 4622 3740 5306
rect 3700 4616 3752 4622
rect 3896 4570 3924 7210
rect 3988 7206 4016 7822
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6798 4016 7142
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4080 6322 4108 8298
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7274 4200 7890
rect 4264 7410 4292 8502
rect 4338 8188 4646 8208
rect 4338 8186 4344 8188
rect 4400 8186 4424 8188
rect 4480 8186 4504 8188
rect 4560 8186 4584 8188
rect 4640 8186 4646 8188
rect 4400 8134 4402 8186
rect 4582 8134 4584 8186
rect 4338 8132 4344 8134
rect 4400 8132 4424 8134
rect 4480 8132 4504 8134
rect 4560 8132 4584 8134
rect 4640 8132 4646 8134
rect 4338 8112 4646 8132
rect 4724 7410 4752 8570
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5000 8022 5028 8434
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6662 4200 7210
rect 4338 7100 4646 7120
rect 4338 7098 4344 7100
rect 4400 7098 4424 7100
rect 4480 7098 4504 7100
rect 4560 7098 4584 7100
rect 4640 7098 4646 7100
rect 4400 7046 4402 7098
rect 4582 7046 4584 7098
rect 4338 7044 4344 7046
rect 4400 7044 4424 7046
rect 4480 7044 4504 7046
rect 4560 7044 4584 7046
rect 4640 7044 4646 7046
rect 4338 7024 4646 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4264 6866 4292 6938
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6390 4660 6598
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4908 6322 4936 7278
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5234 4200 6054
rect 4338 6012 4646 6032
rect 4338 6010 4344 6012
rect 4400 6010 4424 6012
rect 4480 6010 4504 6012
rect 4560 6010 4584 6012
rect 4640 6010 4646 6012
rect 4400 5958 4402 6010
rect 4582 5958 4584 6010
rect 4338 5956 4344 5958
rect 4400 5956 4424 5958
rect 4480 5956 4504 5958
rect 4560 5956 4584 5958
rect 4640 5956 4646 5958
rect 4338 5936 4646 5956
rect 4724 5642 4752 6258
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5710 4844 6190
rect 5000 5914 5028 6258
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4338 4924 4646 4944
rect 4338 4922 4344 4924
rect 4400 4922 4424 4924
rect 4480 4922 4504 4924
rect 4560 4922 4584 4924
rect 4640 4922 4646 4924
rect 4400 4870 4402 4922
rect 4582 4870 4584 4922
rect 4338 4868 4344 4870
rect 4400 4868 4424 4870
rect 4480 4868 4504 4870
rect 4560 4868 4584 4870
rect 4640 4868 4646 4870
rect 4338 4848 4646 4868
rect 4724 4622 4752 5578
rect 4712 4616 4764 4622
rect 3700 4558 3752 4564
rect 3804 4542 4016 4570
rect 4712 4558 4764 4564
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3641 3280 4082
rect 3712 3738 3740 4150
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3238 3632 3294 3641
rect 3238 3567 3294 3576
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 3712 3058 3740 3674
rect 3804 3126 3832 4542
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 3942 3924 4422
rect 3988 4128 4016 4542
rect 4160 4140 4212 4146
rect 3988 4100 4160 4128
rect 4160 4082 4212 4088
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3988 3534 4016 3946
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3976 3392 4028 3398
rect 3974 3360 3976 3369
rect 4028 3360 4030 3369
rect 3974 3295 4030 3304
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 2976 800 3004 2314
rect 3528 800 3556 2858
rect 4080 800 4108 3878
rect 4264 3670 4292 4014
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4338 3836 4646 3856
rect 4338 3834 4344 3836
rect 4400 3834 4424 3836
rect 4480 3834 4504 3836
rect 4560 3834 4584 3836
rect 4640 3834 4646 3836
rect 4400 3782 4402 3834
rect 4582 3782 4584 3834
rect 4338 3780 4344 3782
rect 4400 3780 4424 3782
rect 4480 3780 4504 3782
rect 4560 3780 4584 3782
rect 4640 3780 4646 3782
rect 4338 3760 4646 3780
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4526 3632 4582 3641
rect 4356 3466 4384 3606
rect 4526 3567 4582 3576
rect 4540 3534 4568 3567
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4172 2582 4200 3402
rect 4540 3398 4568 3470
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4338 2748 4646 2768
rect 4338 2746 4344 2748
rect 4400 2746 4424 2748
rect 4480 2746 4504 2748
rect 4560 2746 4584 2748
rect 4640 2746 4646 2748
rect 4400 2694 4402 2746
rect 4582 2694 4584 2746
rect 4338 2692 4344 2694
rect 4400 2692 4424 2694
rect 4480 2692 4504 2694
rect 4560 2692 4584 2694
rect 4640 2692 4646 2694
rect 4338 2672 4646 2692
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 4356 2106 4384 2246
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 4724 1442 4752 3946
rect 4816 3398 4844 5646
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 4908 4826 4936 5578
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5092 4570 5120 9998
rect 5276 9674 5304 11648
rect 5356 11630 5408 11636
rect 5460 10062 5488 12158
rect 5644 11150 5672 12718
rect 5828 11150 5856 12854
rect 6012 12238 6040 15030
rect 6104 12782 6132 15150
rect 6182 14784 6238 14793
rect 6182 14719 6238 14728
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6196 12374 6224 14719
rect 6288 14618 6316 16186
rect 6380 16182 6408 16934
rect 6368 16176 6420 16182
rect 6368 16118 6420 16124
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6472 13462 6500 19306
rect 6564 18426 6592 21490
rect 6932 20602 6960 21966
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6642 20496 6698 20505
rect 6642 20431 6644 20440
rect 6696 20431 6698 20440
rect 6644 20402 6696 20408
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18970 6684 19314
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6748 18902 6776 19722
rect 6840 19378 6868 20198
rect 7024 19922 7052 20334
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6736 18760 6788 18766
rect 6734 18728 6736 18737
rect 6788 18728 6790 18737
rect 6734 18663 6790 18672
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6564 17882 6592 18158
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6656 17678 6684 18226
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6748 17678 6776 18090
rect 6644 17672 6696 17678
rect 6564 17632 6644 17660
rect 6564 17338 6592 17632
rect 6644 17614 6696 17620
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6840 17202 6868 17546
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6840 16046 6868 16662
rect 6828 16040 6880 16046
rect 6550 16008 6606 16017
rect 6828 15982 6880 15988
rect 6550 15943 6606 15952
rect 6564 15638 6592 15943
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6564 12986 6592 15302
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 13326 6684 14010
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6000 12232 6052 12238
rect 5998 12200 6000 12209
rect 6052 12200 6054 12209
rect 5920 12158 5998 12186
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5644 10674 5672 10746
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5448 10056 5500 10062
rect 5184 9646 5304 9674
rect 5368 10016 5448 10044
rect 5184 9042 5212 9646
rect 5368 9586 5396 10016
rect 5448 9998 5500 10004
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5460 9722 5488 9862
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5184 8430 5212 8978
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5184 6746 5212 8366
rect 5276 7886 5304 8978
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8634 5396 8774
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5460 8022 5488 9658
rect 5644 9586 5672 9998
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 8090 5580 8502
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5644 7954 5672 9318
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7478 5304 7822
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 7002 5396 7346
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5356 6792 5408 6798
rect 5184 6718 5304 6746
rect 5356 6734 5408 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6458 5212 6598
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5276 6202 5304 6718
rect 5368 6633 5396 6734
rect 5354 6624 5410 6633
rect 5354 6559 5410 6568
rect 5184 6174 5304 6202
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5184 5846 5212 6174
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4908 4542 5120 4570
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4908 2990 4936 4542
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 2990 5028 4082
rect 5092 4078 5120 4422
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5184 3602 5212 5782
rect 5276 5778 5304 5850
rect 5368 5778 5396 6190
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5276 5234 5304 5714
rect 5368 5574 5396 5714
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5234 5396 5510
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 3670 5396 4558
rect 5460 4010 5488 7686
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 4282 5580 6598
rect 5644 4622 5672 7890
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3194 5396 3334
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5552 3058 5580 3674
rect 5644 3534 5672 4558
rect 5736 3602 5764 11018
rect 5828 4758 5856 11086
rect 5920 8974 5948 12158
rect 5998 12135 6054 12144
rect 6196 11694 6224 12310
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6550 12200 6606 12209
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6288 11354 6316 12174
rect 6550 12135 6606 12144
rect 6564 11762 6592 12135
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6288 11082 6316 11290
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6642 10568 6698 10577
rect 6642 10503 6698 10512
rect 6656 10470 6684 10503
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 6012 8906 6040 9386
rect 6104 9178 6132 9522
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6196 9042 6224 9318
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5920 4214 5948 7346
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6798 6040 7142
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6104 6186 6132 8910
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6196 4622 6224 7686
rect 6288 6202 6316 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6380 8430 6408 9658
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 7410 6408 8366
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6472 6458 6500 10134
rect 6656 8294 6684 10406
rect 6748 9058 6776 15846
rect 6932 15552 6960 18566
rect 7024 18426 7052 19382
rect 7116 19174 7144 22066
rect 7576 22030 7604 23911
rect 8312 22030 8340 23911
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 7727 21788 8035 21808
rect 7727 21786 7733 21788
rect 7789 21786 7813 21788
rect 7869 21786 7893 21788
rect 7949 21786 7973 21788
rect 8029 21786 8035 21788
rect 7789 21734 7791 21786
rect 7971 21734 7973 21786
rect 7727 21732 7733 21734
rect 7789 21732 7813 21734
rect 7869 21732 7893 21734
rect 7949 21732 7973 21734
rect 8029 21732 8035 21734
rect 7727 21712 8035 21732
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7208 19922 7236 21014
rect 7378 20632 7434 20641
rect 7378 20567 7434 20576
rect 7392 20534 7420 20567
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7380 20528 7432 20534
rect 7380 20470 7432 20476
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7208 18952 7236 19858
rect 7300 19854 7328 20470
rect 7484 20262 7512 21422
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7288 19848 7340 19854
rect 7576 19825 7604 21354
rect 8036 21146 8064 21422
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 20466 7696 20742
rect 7727 20700 8035 20720
rect 7727 20698 7733 20700
rect 7789 20698 7813 20700
rect 7869 20698 7893 20700
rect 7949 20698 7973 20700
rect 8029 20698 8035 20700
rect 7789 20646 7791 20698
rect 7971 20646 7973 20698
rect 7727 20644 7733 20646
rect 7789 20644 7813 20646
rect 7869 20644 7893 20646
rect 7949 20644 7973 20646
rect 8029 20644 8035 20646
rect 7727 20624 8035 20644
rect 8128 20602 8156 20810
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7668 19922 7696 20198
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7760 19854 7788 20334
rect 7852 19854 7880 20402
rect 8128 19922 8156 20538
rect 8220 20466 8248 20878
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8220 19990 8248 20402
rect 8312 20330 8340 21490
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 7748 19848 7800 19854
rect 7288 19790 7340 19796
rect 7562 19816 7618 19825
rect 7300 19378 7328 19790
rect 7748 19790 7800 19796
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7562 19751 7618 19760
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 7727 19612 8035 19632
rect 7727 19610 7733 19612
rect 7789 19610 7813 19612
rect 7869 19610 7893 19612
rect 7949 19610 7973 19612
rect 8029 19610 8035 19612
rect 7789 19558 7791 19610
rect 7971 19558 7973 19610
rect 7727 19556 7733 19558
rect 7789 19556 7813 19558
rect 7869 19556 7893 19558
rect 7949 19556 7973 19558
rect 8029 19556 8035 19558
rect 7727 19536 8035 19556
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7208 18924 7420 18952
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7196 18760 7248 18766
rect 7194 18728 7196 18737
rect 7248 18728 7250 18737
rect 7194 18663 7250 18672
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7300 18358 7328 18770
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 17338 7052 18022
rect 7208 17678 7236 18294
rect 7392 18204 7420 18924
rect 7300 18176 7420 18204
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7024 16590 7052 17138
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7116 16250 7144 16934
rect 7208 16794 7236 17614
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7208 16454 7236 16730
rect 7300 16590 7328 18176
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7392 16794 7420 17070
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7288 16584 7340 16590
rect 7286 16552 7288 16561
rect 7340 16552 7342 16561
rect 7392 16522 7420 16730
rect 7484 16590 7512 17070
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7286 16487 7342 16496
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7576 15570 7604 17614
rect 7668 16454 7696 19314
rect 7727 18524 8035 18544
rect 7727 18522 7733 18524
rect 7789 18522 7813 18524
rect 7869 18522 7893 18524
rect 7949 18522 7973 18524
rect 8029 18522 8035 18524
rect 7789 18470 7791 18522
rect 7971 18470 7973 18522
rect 7727 18468 7733 18470
rect 7789 18468 7813 18470
rect 7869 18468 7893 18470
rect 7949 18468 7973 18470
rect 8029 18468 8035 18470
rect 7727 18448 8035 18468
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 17814 7880 18226
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7727 17436 8035 17456
rect 7727 17434 7733 17436
rect 7789 17434 7813 17436
rect 7869 17434 7893 17436
rect 7949 17434 7973 17436
rect 8029 17434 8035 17436
rect 7789 17382 7791 17434
rect 7971 17382 7973 17434
rect 7727 17380 7733 17382
rect 7789 17380 7813 17382
rect 7869 17380 7893 17382
rect 7949 17380 7973 17382
rect 8029 17380 8035 17382
rect 7727 17360 8035 17380
rect 8128 16522 8156 19722
rect 8220 16776 8248 19790
rect 8300 18284 8352 18290
rect 8404 18272 8432 20470
rect 8496 19786 8524 20946
rect 8680 20602 8708 21286
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8758 20496 8814 20505
rect 8668 20460 8720 20466
rect 8758 20431 8760 20440
rect 8668 20402 8720 20408
rect 8812 20431 8814 20440
rect 8760 20402 8812 20408
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8352 18244 8432 18272
rect 8300 18226 8352 18232
rect 8312 17270 8340 18226
rect 8496 17678 8524 19382
rect 8588 18290 8616 20198
rect 8680 20058 8708 20402
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8680 19514 8708 19790
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8772 19378 8800 20402
rect 8864 20058 8892 23911
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8484 17672 8536 17678
rect 8482 17640 8484 17649
rect 8536 17640 8538 17649
rect 8482 17575 8538 17584
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8220 16748 8340 16776
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7727 16348 8035 16368
rect 7727 16346 7733 16348
rect 7789 16346 7813 16348
rect 7869 16346 7893 16348
rect 7949 16346 7973 16348
rect 8029 16346 8035 16348
rect 7789 16294 7791 16346
rect 7971 16294 7973 16346
rect 7727 16292 7733 16294
rect 7789 16292 7813 16294
rect 7869 16292 7893 16294
rect 7949 16292 7973 16294
rect 8029 16292 8035 16294
rect 7727 16272 8035 16292
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7104 15564 7156 15570
rect 6932 15524 7052 15552
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14414 6868 14758
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 12730 6868 13806
rect 6932 13802 6960 14894
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6840 12702 6960 12730
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12238 6868 12582
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11694 6868 12174
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 10606 6868 11630
rect 6932 11286 6960 12702
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10674 6960 10950
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 9722 6868 10406
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9722 6960 10066
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6840 9382 6868 9658
rect 7024 9586 7052 15524
rect 7564 15564 7616 15570
rect 7104 15506 7156 15512
rect 7484 15524 7564 15552
rect 7116 11830 7144 15506
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 15094 7420 15438
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7392 14482 7420 15030
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7208 14006 7236 14418
rect 7288 14408 7340 14414
rect 7484 14362 7512 15524
rect 7564 15506 7616 15512
rect 7668 15162 7696 16050
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7727 15260 8035 15280
rect 7727 15258 7733 15260
rect 7789 15258 7813 15260
rect 7869 15258 7893 15260
rect 7949 15258 7973 15260
rect 8029 15258 8035 15260
rect 7789 15206 7791 15258
rect 7971 15206 7973 15258
rect 7727 15204 7733 15206
rect 7789 15204 7813 15206
rect 7869 15204 7893 15206
rect 7949 15204 7973 15206
rect 8029 15204 8035 15206
rect 7727 15184 8035 15204
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7288 14350 7340 14356
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7208 12646 7236 13942
rect 7300 13258 7328 14350
rect 7392 14334 7512 14362
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7300 12442 7328 13194
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7116 9654 7144 11766
rect 7208 11354 7236 12174
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 7208 9194 7236 11086
rect 7300 10266 7328 12378
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7024 9166 7236 9194
rect 6748 9030 6868 9058
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8634 6776 8910
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6564 6798 6592 7414
rect 6656 7188 6684 8230
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6748 7546 6776 7890
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6736 7200 6788 7206
rect 6656 7160 6736 7188
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6288 6174 6408 6202
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5710 6316 6054
rect 6380 5817 6408 6174
rect 6366 5808 6422 5817
rect 6366 5743 6422 5752
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 5370 6408 5510
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6472 5114 6500 6394
rect 6380 5086 6500 5114
rect 6380 4826 6408 5086
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 6196 4146 6224 4558
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6196 3534 6224 4082
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3534 6408 3878
rect 6472 3738 6500 4966
rect 6656 3942 6684 7160
rect 6736 7142 6788 7148
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 4214 6776 6054
rect 6840 4622 6868 9030
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6932 6934 6960 8842
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 7024 6610 7052 9166
rect 7194 9072 7250 9081
rect 7104 9036 7156 9042
rect 7194 9007 7250 9016
rect 7104 8978 7156 8984
rect 7116 6866 7144 8978
rect 7208 8974 7236 9007
rect 7300 8974 7328 10202
rect 7392 10033 7420 14334
rect 7470 14104 7526 14113
rect 7470 14039 7526 14048
rect 7484 13938 7512 14039
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13326 7512 13874
rect 7576 13394 7604 14554
rect 7668 14074 7696 15098
rect 7746 15056 7802 15065
rect 7746 14991 7748 15000
rect 7800 14991 7802 15000
rect 7748 14962 7800 14968
rect 8220 14958 8248 15914
rect 8312 15366 8340 16748
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 7727 14172 8035 14192
rect 7727 14170 7733 14172
rect 7789 14170 7813 14172
rect 7869 14170 7893 14172
rect 7949 14170 7973 14172
rect 8029 14170 8035 14172
rect 7789 14118 7791 14170
rect 7971 14118 7973 14170
rect 7727 14116 7733 14118
rect 7789 14116 7813 14118
rect 7869 14116 7893 14118
rect 7949 14116 7973 14118
rect 8029 14116 8035 14118
rect 7727 14096 8035 14116
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 8128 14006 8156 14826
rect 8404 14822 8432 16118
rect 8496 15858 8524 17478
rect 8588 16980 8616 18226
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8680 17202 8708 17682
rect 8772 17678 8800 18158
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8850 17232 8906 17241
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8668 16992 8720 16998
rect 8588 16952 8668 16980
rect 8668 16934 8720 16940
rect 8496 15830 8616 15858
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7484 12782 7512 12854
rect 7668 12850 7696 13398
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7727 13084 8035 13104
rect 7727 13082 7733 13084
rect 7789 13082 7813 13084
rect 7869 13082 7893 13084
rect 7949 13082 7973 13084
rect 8029 13082 8035 13084
rect 7789 13030 7791 13082
rect 7971 13030 7973 13082
rect 7727 13028 7733 13030
rect 7789 13028 7813 13030
rect 7869 13028 7893 13030
rect 7949 13028 7973 13030
rect 8029 13028 8035 13030
rect 7727 13008 8035 13028
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7472 12776 7524 12782
rect 7524 12736 7604 12764
rect 7472 12718 7524 12724
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7378 10024 7434 10033
rect 7378 9959 7434 9968
rect 7392 9518 7420 9959
rect 7484 9738 7512 12582
rect 7576 12238 7604 12736
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7668 11880 7696 12786
rect 8128 12306 8156 13330
rect 8220 12374 8248 14010
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7727 11996 8035 12016
rect 7727 11994 7733 11996
rect 7789 11994 7813 11996
rect 7869 11994 7893 11996
rect 7949 11994 7973 11996
rect 8029 11994 8035 11996
rect 7789 11942 7791 11994
rect 7971 11942 7973 11994
rect 7727 11940 7733 11942
rect 7789 11940 7813 11942
rect 7869 11940 7893 11942
rect 7949 11940 7973 11942
rect 8029 11940 8035 11942
rect 7727 11920 8035 11940
rect 7668 11852 7788 11880
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7576 10577 7604 11154
rect 7668 11150 7696 11494
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7760 10996 7788 11852
rect 7668 10968 7788 10996
rect 7668 10810 7696 10968
rect 7727 10908 8035 10928
rect 7727 10906 7733 10908
rect 7789 10906 7813 10908
rect 7869 10906 7893 10908
rect 7949 10906 7973 10908
rect 8029 10906 8035 10908
rect 7789 10854 7791 10906
rect 7971 10854 7973 10906
rect 7727 10852 7733 10854
rect 7789 10852 7813 10854
rect 7869 10852 7893 10854
rect 7949 10852 7973 10854
rect 8029 10852 8035 10854
rect 7727 10832 8035 10852
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7668 10674 7696 10746
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7562 10568 7618 10577
rect 7562 10503 7618 10512
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7576 10062 7604 10406
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7484 9710 7604 9738
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7208 7206 7236 8910
rect 7392 7886 7420 9046
rect 7484 8906 7512 9522
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 8498 7512 8842
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7300 7041 7328 7686
rect 7484 7546 7512 8298
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7286 7032 7342 7041
rect 7286 6967 7342 6976
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7024 6582 7144 6610
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7010 6216 7066 6225
rect 6932 6118 6960 6190
rect 7010 6151 7066 6160
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6932 4486 6960 5102
rect 7024 5030 7052 6151
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7116 4593 7144 6582
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7102 4584 7158 4593
rect 7012 4548 7064 4554
rect 7102 4519 7158 4528
rect 7012 4490 7064 4496
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6932 3670 6960 4422
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7024 3534 7052 4490
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 5644 3058 5672 3470
rect 6196 3194 6224 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3194 7052 3334
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 7116 2774 7144 4422
rect 7208 4128 7236 6258
rect 7300 5234 7328 6870
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6458 7420 6734
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7484 6361 7512 7482
rect 7470 6352 7526 6361
rect 7470 6287 7526 6296
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5302 7420 6054
rect 7484 5914 7512 6151
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7484 5234 7512 5646
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7300 4282 7328 4966
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7208 4100 7420 4128
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7300 3534 7328 3946
rect 7392 3534 7420 4100
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7300 2990 7328 3062
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7024 2746 7144 2774
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 4632 1414 4752 1442
rect 4632 800 4660 1414
rect 5368 800 5396 2382
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5920 800 5948 2314
rect 6472 800 6500 2382
rect 7024 800 7052 2746
rect 7576 2038 7604 9710
rect 7668 9042 7696 10406
rect 7852 10266 7880 10610
rect 8128 10470 8156 12242
rect 8220 11014 8248 12310
rect 8312 12209 8340 13806
rect 8404 13802 8432 14758
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8298 12200 8354 12209
rect 8298 12135 8354 12144
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11898 8340 12038
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7727 9820 8035 9840
rect 7727 9818 7733 9820
rect 7789 9818 7813 9820
rect 7869 9818 7893 9820
rect 7949 9818 7973 9820
rect 8029 9818 8035 9820
rect 7789 9766 7791 9818
rect 7971 9766 7973 9818
rect 7727 9764 7733 9766
rect 7789 9764 7813 9766
rect 7869 9764 7893 9766
rect 7949 9764 7973 9766
rect 8029 9764 8035 9766
rect 7727 9744 8035 9764
rect 8128 9625 8156 9998
rect 8114 9616 8170 9625
rect 8114 9551 8170 9560
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7748 8968 7800 8974
rect 7668 8916 7748 8922
rect 7668 8910 7800 8916
rect 7668 8894 7788 8910
rect 7668 8566 7696 8894
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7727 8732 8035 8752
rect 7727 8730 7733 8732
rect 7789 8730 7813 8732
rect 7869 8730 7893 8732
rect 7949 8730 7973 8732
rect 8029 8730 8035 8732
rect 7789 8678 7791 8730
rect 7971 8678 7973 8730
rect 7727 8676 7733 8678
rect 7789 8676 7813 8678
rect 7869 8676 7893 8678
rect 7949 8676 7973 8678
rect 8029 8676 8035 8678
rect 7727 8656 8035 8676
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 8128 8430 8156 8774
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7838 7984 7894 7993
rect 7838 7919 7840 7928
rect 7892 7919 7894 7928
rect 7840 7890 7892 7896
rect 7727 7644 8035 7664
rect 7727 7642 7733 7644
rect 7789 7642 7813 7644
rect 7869 7642 7893 7644
rect 7949 7642 7973 7644
rect 8029 7642 8035 7644
rect 7789 7590 7791 7642
rect 7971 7590 7973 7642
rect 7727 7588 7733 7590
rect 7789 7588 7813 7590
rect 7869 7588 7893 7590
rect 7949 7588 7973 7590
rect 8029 7588 8035 7590
rect 7727 7568 8035 7588
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8128 6934 8156 7278
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7668 5710 7696 6802
rect 8220 6712 8248 10610
rect 8298 10296 8354 10305
rect 8298 10231 8300 10240
rect 8352 10231 8354 10240
rect 8300 10202 8352 10208
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8312 9450 8340 9658
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8298 7440 8354 7449
rect 8298 7375 8300 7384
rect 8352 7375 8354 7384
rect 8300 7346 8352 7352
rect 8312 7002 8340 7346
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8404 6866 8432 13262
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8128 6684 8248 6712
rect 8392 6724 8444 6730
rect 7727 6556 8035 6576
rect 7727 6554 7733 6556
rect 7789 6554 7813 6556
rect 7869 6554 7893 6556
rect 7949 6554 7973 6556
rect 8029 6554 8035 6556
rect 7789 6502 7791 6554
rect 7971 6502 7973 6554
rect 7727 6500 7733 6502
rect 7789 6500 7813 6502
rect 7869 6500 7893 6502
rect 7949 6500 7973 6502
rect 8029 6500 8035 6502
rect 7727 6480 8035 6500
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7668 5098 7696 5510
rect 7727 5468 8035 5488
rect 7727 5466 7733 5468
rect 7789 5466 7813 5468
rect 7869 5466 7893 5468
rect 7949 5466 7973 5468
rect 8029 5466 8035 5468
rect 7789 5414 7791 5466
rect 7971 5414 7973 5466
rect 7727 5412 7733 5414
rect 7789 5412 7813 5414
rect 7869 5412 7893 5414
rect 7949 5412 7973 5414
rect 8029 5412 8035 5414
rect 7727 5392 8035 5412
rect 7748 5228 7800 5234
rect 7800 5188 7880 5216
rect 7748 5170 7800 5176
rect 7852 5098 7880 5188
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4622 7788 4966
rect 7748 4616 7800 4622
rect 7668 4576 7748 4604
rect 7668 3738 7696 4576
rect 7748 4558 7800 4564
rect 7852 4554 7880 5034
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7727 4380 8035 4400
rect 7727 4378 7733 4380
rect 7789 4378 7813 4380
rect 7869 4378 7893 4380
rect 7949 4378 7973 4380
rect 8029 4378 8035 4380
rect 7789 4326 7791 4378
rect 7971 4326 7973 4378
rect 7727 4324 7733 4326
rect 7789 4324 7813 4326
rect 7869 4324 7893 4326
rect 7949 4324 7973 4326
rect 8029 4324 8035 4326
rect 7727 4304 8035 4324
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 8036 3534 8064 4082
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7727 3292 8035 3312
rect 7727 3290 7733 3292
rect 7789 3290 7813 3292
rect 7869 3290 7893 3292
rect 7949 3290 7973 3292
rect 8029 3290 8035 3292
rect 7789 3238 7791 3290
rect 7971 3238 7973 3290
rect 7727 3236 7733 3238
rect 7789 3236 7813 3238
rect 7869 3236 7893 3238
rect 7949 3236 7973 3238
rect 8029 3236 8035 3238
rect 7727 3216 8035 3236
rect 7727 2204 8035 2224
rect 7727 2202 7733 2204
rect 7789 2202 7813 2204
rect 7869 2202 7893 2204
rect 7949 2202 7973 2204
rect 8029 2202 8035 2204
rect 7789 2150 7791 2202
rect 7971 2150 7973 2202
rect 7727 2148 7733 2150
rect 7789 2148 7813 2150
rect 7869 2148 7893 2150
rect 7949 2148 7973 2150
rect 8029 2148 8035 2150
rect 7727 2128 8035 2148
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7760 870 7880 898
rect 7760 800 7788 870
rect 18 0 74 800
rect 570 0 626 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3514 0 3570 800
rect 4066 0 4122 800
rect 4618 0 4674 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7746 0 7802 800
rect 7852 762 7880 870
rect 8128 762 8156 6684
rect 8392 6666 8444 6672
rect 8404 6322 8432 6666
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 2922 8248 4490
rect 8312 4214 8340 6054
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3194 8340 3878
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 3074 8432 3130
rect 8312 3058 8432 3074
rect 8300 3052 8432 3058
rect 8352 3046 8432 3052
rect 8300 2994 8352 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8496 2582 8524 15642
rect 8588 13462 8616 15830
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8680 11898 8708 16934
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11082 8616 11630
rect 8772 11286 8800 17206
rect 8850 17167 8906 17176
rect 8864 17134 8892 17167
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16726 8892 17070
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14414 8892 14758
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 14006 8892 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8864 13394 8892 13942
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 13025 8892 13126
rect 8850 13016 8906 13025
rect 8850 12951 8906 12960
rect 8864 12850 8892 12951
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8956 12434 8984 21830
rect 9416 21690 9444 23911
rect 9968 22030 9996 23911
rect 10704 23882 10732 23911
rect 10796 23882 10824 23990
rect 10704 23854 10824 23882
rect 10980 22094 11008 23990
rect 11242 23911 11298 24711
rect 11348 23990 11560 24018
rect 11256 23882 11284 23911
rect 11348 23882 11376 23990
rect 11256 23854 11376 23882
rect 11116 22332 11424 22352
rect 11116 22330 11122 22332
rect 11178 22330 11202 22332
rect 11258 22330 11282 22332
rect 11338 22330 11362 22332
rect 11418 22330 11424 22332
rect 11178 22278 11180 22330
rect 11360 22278 11362 22330
rect 11116 22276 11122 22278
rect 11178 22276 11202 22278
rect 11258 22276 11282 22278
rect 11338 22276 11362 22278
rect 11418 22276 11424 22278
rect 11116 22256 11424 22276
rect 11152 22094 11204 22098
rect 10980 22092 11204 22094
rect 10980 22066 11152 22092
rect 11152 22034 11204 22040
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10600 22024 10652 22030
rect 10876 22024 10928 22030
rect 10600 21966 10652 21972
rect 10704 21984 10876 22012
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 9312 21616 9364 21622
rect 9312 21558 9364 21564
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9140 20806 9168 21354
rect 9232 20942 9260 21422
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 9324 19854 9352 21558
rect 10244 21554 10272 21626
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10060 21457 10088 21490
rect 10046 21448 10102 21457
rect 10046 21383 10102 21392
rect 10244 21406 10456 21434
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9588 21004 9640 21010
rect 9772 21004 9824 21010
rect 9640 20964 9772 20992
rect 9588 20946 9640 20952
rect 9772 20946 9824 20952
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9600 19854 9628 20266
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 9048 18970 9076 19722
rect 9324 19417 9352 19790
rect 9310 19408 9366 19417
rect 9128 19372 9180 19378
rect 9310 19343 9312 19352
rect 9128 19314 9180 19320
rect 9364 19343 9366 19352
rect 9312 19314 9364 19320
rect 9140 19258 9168 19314
rect 9140 19230 9352 19258
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9048 17814 9076 18702
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 18290 9168 18566
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9140 17746 9168 18226
rect 9232 17882 9260 18226
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9036 17672 9088 17678
rect 9324 17660 9352 19230
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9508 17678 9536 17818
rect 9496 17672 9548 17678
rect 9324 17632 9444 17660
rect 9036 17614 9088 17620
rect 9048 15706 9076 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9232 15502 9260 16730
rect 9324 16658 9352 17478
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9324 16561 9352 16594
rect 9310 16552 9366 16561
rect 9310 16487 9366 16496
rect 9416 15570 9444 17632
rect 9496 17614 9548 17620
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 13734 9076 15302
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9232 14618 9260 15030
rect 9310 14920 9366 14929
rect 9310 14855 9366 14864
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9324 14414 9352 14855
rect 9508 14657 9536 17614
rect 9600 16998 9628 19790
rect 9692 19718 9720 20470
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9784 19553 9812 20538
rect 9876 20466 9904 21082
rect 9968 20482 9996 21286
rect 10138 21040 10194 21049
rect 10138 20975 10194 20984
rect 10152 20942 10180 20975
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10048 20800 10100 20806
rect 10046 20768 10048 20777
rect 10100 20768 10102 20777
rect 10046 20703 10102 20712
rect 10244 20602 10272 21406
rect 10428 21350 10456 21406
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10336 20942 10364 21286
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10428 20602 10456 20946
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 9864 20460 9916 20466
rect 9968 20454 10364 20482
rect 9864 20402 9916 20408
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 19922 9996 20198
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9770 19544 9826 19553
rect 9876 19514 9904 19654
rect 9770 19479 9826 19488
rect 9864 19508 9916 19514
rect 9784 19378 9812 19479
rect 9864 19450 9916 19456
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9784 17338 9812 18158
rect 9968 17814 9996 19314
rect 10060 18222 10088 19858
rect 10244 19378 10272 20266
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10152 18698 10180 19314
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18766 10272 19110
rect 10336 18902 10364 20454
rect 10324 18896 10376 18902
rect 10376 18856 10456 18884
rect 10324 18838 10376 18844
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9692 15706 9720 16458
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9494 14648 9550 14657
rect 9494 14583 9550 14592
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9218 14104 9274 14113
rect 9218 14039 9274 14048
rect 9494 14104 9550 14113
rect 9494 14039 9550 14048
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12850 9076 13126
rect 9140 12918 9168 13330
rect 9232 13190 9260 14039
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9128 12640 9180 12646
rect 9126 12608 9128 12617
rect 9180 12608 9182 12617
rect 9126 12543 9182 12552
rect 8864 12406 8984 12434
rect 9126 12472 9182 12481
rect 9126 12407 9182 12416
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8680 10470 8708 10746
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8588 7886 8616 9590
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 8634 8708 9522
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8772 8498 8800 8570
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 5778 8616 7822
rect 8864 7818 8892 12406
rect 9140 11626 9168 12407
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 10742 8984 11494
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8956 10266 8984 10474
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9761 8984 9862
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8956 8974 8984 9114
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8956 7698 8984 8910
rect 9048 7886 9076 9454
rect 9140 8090 9168 11086
rect 9232 10606 9260 13126
rect 9324 11762 9352 13466
rect 9416 13462 9444 13670
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9508 13326 9536 14039
rect 9600 13734 9628 15506
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14521 9720 14758
rect 9678 14512 9734 14521
rect 9678 14447 9734 14456
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9784 12986 9812 16934
rect 10060 16266 10088 18158
rect 10152 17678 10180 18634
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18426 10364 18566
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10230 17776 10286 17785
rect 10230 17711 10286 17720
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10244 17610 10272 17711
rect 10336 17678 10364 18226
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10230 16688 10286 16697
rect 10230 16623 10232 16632
rect 10284 16623 10286 16632
rect 10232 16594 10284 16600
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10060 16238 10180 16266
rect 10244 16250 10272 16390
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 10060 15910 10088 16118
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9876 15502 9904 15846
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 15162 9996 15438
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 14278 9904 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9968 14074 9996 14894
rect 10060 14618 10088 15574
rect 10152 15094 10180 16238
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10230 16008 10286 16017
rect 10230 15943 10286 15952
rect 10244 15910 10272 15943
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10140 15088 10192 15094
rect 10192 15048 10272 15076
rect 10140 15030 10192 15036
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9954 13968 10010 13977
rect 9954 13903 10010 13912
rect 9968 13734 9996 13903
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 10060 13530 10088 14554
rect 10152 13938 10180 14758
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 13394 10088 13466
rect 10244 13462 10272 15048
rect 10140 13456 10192 13462
rect 10138 13424 10140 13433
rect 10232 13456 10284 13462
rect 10192 13424 10194 13433
rect 10048 13388 10100 13394
rect 10232 13398 10284 13404
rect 10138 13359 10194 13368
rect 10048 13330 10100 13336
rect 10244 13274 10272 13398
rect 10152 13246 10272 13274
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9402 12608 9458 12617
rect 9402 12543 9458 12552
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11354 9352 11698
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9220 10464 9272 10470
rect 9416 10418 9444 12543
rect 9508 12442 9536 12650
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9494 12336 9550 12345
rect 9494 12271 9550 12280
rect 9220 10406 9272 10412
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8864 7670 8984 7698
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 2990 8616 5714
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8772 2922 8800 7346
rect 8864 4706 8892 7670
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8956 4842 8984 6734
rect 9048 6322 9076 7822
rect 9126 6896 9182 6905
rect 9126 6831 9182 6840
rect 9140 6662 9168 6831
rect 9232 6798 9260 10406
rect 9324 10390 9444 10418
rect 9324 8294 9352 10390
rect 9508 10266 9536 12271
rect 9600 11558 9628 12786
rect 9862 12744 9918 12753
rect 9862 12679 9918 12688
rect 9876 12646 9904 12679
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 10152 11830 10180 13246
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10244 12986 10272 13126
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10336 12866 10364 17614
rect 10428 16658 10456 18856
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10428 15502 10456 16050
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14822 10456 15438
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 12986 10456 13806
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10244 12838 10364 12866
rect 10428 12850 10456 12922
rect 10416 12844 10468 12850
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9784 11150 9812 11766
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9232 5658 9260 6734
rect 9324 5914 9352 7142
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9140 5630 9260 5658
rect 9034 5536 9090 5545
rect 9034 5471 9090 5480
rect 9048 5370 9076 5471
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9140 5234 9168 5630
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 5370 9260 5510
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9324 5273 9352 5714
rect 9310 5264 9366 5273
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9220 5228 9272 5234
rect 9310 5199 9366 5208
rect 9220 5170 9272 5176
rect 9232 4865 9260 5170
rect 9218 4856 9274 4865
rect 8956 4814 9168 4842
rect 9036 4752 9088 4758
rect 8864 4678 8984 4706
rect 9036 4694 9088 4700
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 800 8340 2314
rect 8864 800 8892 4490
rect 8956 2514 8984 4678
rect 9048 4282 9076 4694
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9048 3942 9076 4218
rect 9140 3942 9168 4814
rect 9416 4826 9444 10202
rect 9600 10130 9628 11018
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9494 10024 9550 10033
rect 9494 9959 9550 9968
rect 9508 9926 9536 9959
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9494 9752 9550 9761
rect 9494 9687 9496 9696
rect 9548 9687 9550 9696
rect 9496 9658 9548 9664
rect 9508 9178 9536 9658
rect 9600 9450 9628 10066
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9508 6458 9536 8502
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9600 7546 9628 7822
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6866 9628 7346
rect 9692 7342 9720 7822
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9600 5846 9628 6666
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5545 9536 5578
rect 9494 5536 9550 5545
rect 9494 5471 9550 5480
rect 9600 5409 9628 5646
rect 9586 5400 9642 5409
rect 9586 5335 9642 5344
rect 9692 5302 9720 5782
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9586 5128 9642 5137
rect 9586 5063 9588 5072
rect 9640 5063 9642 5072
rect 9588 5034 9640 5040
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9586 4856 9642 4865
rect 9218 4791 9274 4800
rect 9404 4820 9456 4826
rect 9586 4791 9588 4800
rect 9404 4762 9456 4768
rect 9640 4791 9642 4800
rect 9588 4762 9640 4768
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4282 9536 4626
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4486 9628 4558
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9048 3058 9076 3878
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3058 9352 3470
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9324 2650 9352 2994
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9416 800 9444 3946
rect 9600 3194 9628 4422
rect 9692 4282 9720 4966
rect 9784 4672 9812 7958
rect 9876 6730 9904 10474
rect 9954 10296 10010 10305
rect 10060 10266 10088 10610
rect 9954 10231 10010 10240
rect 10048 10260 10100 10266
rect 9968 8566 9996 10231
rect 10048 10202 10100 10208
rect 10060 9722 10088 10202
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 10060 8480 10088 9658
rect 10152 8974 10180 9862
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10060 8452 10180 8480
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7585 9996 8026
rect 9954 7576 10010 7585
rect 9954 7511 10010 7520
rect 9968 7410 9996 7511
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9876 5302 9904 6326
rect 9968 5778 9996 6394
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9968 5166 9996 5510
rect 9864 5160 9916 5166
rect 9862 5128 9864 5137
rect 9956 5160 10008 5166
rect 9916 5128 9918 5137
rect 9956 5102 10008 5108
rect 9862 5063 9918 5072
rect 10060 4690 10088 8298
rect 10152 8022 10180 8452
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7546 10180 7958
rect 10244 7954 10272 12838
rect 10416 12786 10468 12792
rect 10322 12200 10378 12209
rect 10322 12135 10378 12144
rect 10336 11354 10364 12135
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10428 10538 10456 11630
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10414 10296 10470 10305
rect 10414 10231 10416 10240
rect 10468 10231 10470 10240
rect 10416 10202 10468 10208
rect 10520 9625 10548 21830
rect 10612 20466 10640 21966
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10704 20398 10732 21984
rect 10876 21966 10928 21972
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10888 21146 10916 21830
rect 11532 21690 11560 23990
rect 11794 23911 11850 24711
rect 12346 23911 12402 24711
rect 12636 23990 13032 24018
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11428 21616 11480 21622
rect 11480 21564 11652 21570
rect 11428 21558 11652 21564
rect 11440 21542 11652 21558
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11532 21350 11560 21422
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11116 21244 11424 21264
rect 11116 21242 11122 21244
rect 11178 21242 11202 21244
rect 11258 21242 11282 21244
rect 11338 21242 11362 21244
rect 11418 21242 11424 21244
rect 11178 21190 11180 21242
rect 11360 21190 11362 21242
rect 11116 21188 11122 21190
rect 11178 21188 11202 21190
rect 11258 21188 11282 21190
rect 11338 21188 11362 21190
rect 11418 21188 11424 21190
rect 11116 21168 11424 21188
rect 11624 21146 11652 21542
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11058 21040 11114 21049
rect 10784 21004 10836 21010
rect 11058 20975 11060 20984
rect 10784 20946 10836 20952
rect 11112 20975 11114 20984
rect 11060 20946 11112 20952
rect 10796 20913 10824 20946
rect 10782 20904 10838 20913
rect 10782 20839 10838 20848
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10612 18358 10640 19314
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10704 18290 10732 20334
rect 10796 19922 10824 20839
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10888 19786 10916 20538
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10980 19310 11008 20198
rect 11116 20156 11424 20176
rect 11116 20154 11122 20156
rect 11178 20154 11202 20156
rect 11258 20154 11282 20156
rect 11338 20154 11362 20156
rect 11418 20154 11424 20156
rect 11178 20102 11180 20154
rect 11360 20102 11362 20154
rect 11116 20100 11122 20102
rect 11178 20100 11202 20102
rect 11258 20100 11282 20102
rect 11338 20100 11362 20102
rect 11418 20100 11424 20102
rect 11116 20080 11424 20100
rect 11532 20097 11560 20538
rect 11624 20466 11652 20742
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11518 20088 11574 20097
rect 11518 20023 11574 20032
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11532 19310 11560 19926
rect 11716 19530 11744 21966
rect 11808 19990 11836 23911
rect 12360 22012 12388 23911
rect 12440 22024 12492 22030
rect 12360 21984 12440 22012
rect 12440 21966 12492 21972
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11992 20942 12020 21286
rect 12070 21040 12126 21049
rect 12070 20975 12126 20984
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11992 20466 12020 20878
rect 12084 20806 12112 20975
rect 12072 20800 12124 20806
rect 12070 20768 12072 20777
rect 12124 20768 12126 20777
rect 12070 20703 12126 20712
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11992 19718 12020 20402
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11624 19502 11744 19530
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11116 19068 11424 19088
rect 11116 19066 11122 19068
rect 11178 19066 11202 19068
rect 11258 19066 11282 19068
rect 11338 19066 11362 19068
rect 11418 19066 11424 19068
rect 11178 19014 11180 19066
rect 11360 19014 11362 19066
rect 11116 19012 11122 19014
rect 11178 19012 11202 19014
rect 11258 19012 11282 19014
rect 11338 19012 11362 19014
rect 11418 19012 11424 19014
rect 11116 18992 11424 19012
rect 11532 18902 11560 19246
rect 11520 18896 11572 18902
rect 10782 18864 10838 18873
rect 11520 18838 11572 18844
rect 10782 18799 10784 18808
rect 10836 18799 10838 18808
rect 10784 18770 10836 18776
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10704 17678 10732 17818
rect 10692 17672 10744 17678
rect 10744 17632 10824 17660
rect 10692 17614 10744 17620
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 17202 10640 17546
rect 10796 17241 10824 17632
rect 10782 17232 10838 17241
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10692 17196 10744 17202
rect 10888 17202 10916 18702
rect 11532 18630 11560 18838
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11116 17980 11424 18000
rect 11116 17978 11122 17980
rect 11178 17978 11202 17980
rect 11258 17978 11282 17980
rect 11338 17978 11362 17980
rect 11418 17978 11424 17980
rect 11178 17926 11180 17978
rect 11360 17926 11362 17978
rect 11116 17924 11122 17926
rect 11178 17924 11202 17926
rect 11258 17924 11282 17926
rect 11338 17924 11362 17926
rect 11418 17924 11424 17926
rect 11116 17904 11424 17924
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11518 17640 11574 17649
rect 11348 17338 11376 17614
rect 11518 17575 11574 17584
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 10782 17167 10838 17176
rect 10876 17196 10928 17202
rect 10692 17138 10744 17144
rect 10876 17138 10928 17144
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 15094 10640 15506
rect 10704 15162 10732 17138
rect 11532 16998 11560 17575
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 10796 16046 10824 16934
rect 11116 16892 11424 16912
rect 11116 16890 11122 16892
rect 11178 16890 11202 16892
rect 11258 16890 11282 16892
rect 11338 16890 11362 16892
rect 11418 16890 11424 16892
rect 11178 16838 11180 16890
rect 11360 16838 11362 16890
rect 11116 16836 11122 16838
rect 11178 16836 11202 16838
rect 11258 16836 11282 16838
rect 11338 16836 11362 16838
rect 11418 16836 11424 16838
rect 11116 16816 11424 16836
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10784 15428 10836 15434
rect 10836 15388 10916 15416
rect 10784 15370 10836 15376
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14929 10732 14962
rect 10690 14920 10746 14929
rect 10690 14855 10746 14864
rect 10598 14512 10654 14521
rect 10704 14482 10732 14855
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10598 14447 10654 14456
rect 10692 14476 10744 14482
rect 10612 14414 10640 14447
rect 10692 14418 10744 14424
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10704 13938 10732 14214
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10612 13172 10640 13874
rect 10796 13870 10824 14486
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10796 13462 10824 13670
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10692 13184 10744 13190
rect 10612 13144 10692 13172
rect 10692 13126 10744 13132
rect 10704 12918 10732 13126
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10704 12782 10732 12854
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10704 11354 10732 12174
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10704 10674 10732 11290
rect 10796 11150 10824 12174
rect 10888 12102 10916 15388
rect 10980 14793 11008 16390
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11116 15804 11424 15824
rect 11116 15802 11122 15804
rect 11178 15802 11202 15804
rect 11258 15802 11282 15804
rect 11338 15802 11362 15804
rect 11418 15802 11424 15804
rect 11178 15750 11180 15802
rect 11360 15750 11362 15802
rect 11116 15748 11122 15750
rect 11178 15748 11202 15750
rect 11258 15748 11282 15750
rect 11338 15748 11362 15750
rect 11418 15748 11424 15750
rect 11116 15728 11424 15748
rect 11532 15688 11560 15982
rect 11348 15660 11560 15688
rect 11348 15434 11376 15660
rect 11624 15552 11652 19502
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11886 19408 11942 19417
rect 11716 18290 11744 19382
rect 11886 19343 11942 19352
rect 11980 19372 12032 19378
rect 11900 18329 11928 19343
rect 11980 19314 12032 19320
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11992 18970 12020 19314
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11886 18320 11942 18329
rect 11704 18284 11756 18290
rect 11992 18290 12020 18906
rect 12084 18834 12112 19314
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11886 18255 11942 18264
rect 11980 18284 12032 18290
rect 11704 18226 11756 18232
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16590 11744 17138
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11900 16402 11928 18255
rect 11980 18226 12032 18232
rect 11992 17678 12020 18226
rect 12084 18154 12112 18634
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12084 17882 12112 18090
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11978 17368 12034 17377
rect 11978 17303 12034 17312
rect 11992 17270 12020 17303
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 16658 12112 17070
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11978 16552 12034 16561
rect 11978 16487 12034 16496
rect 11992 16454 12020 16487
rect 11532 15524 11652 15552
rect 11716 16374 11928 16402
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11532 15026 11560 15524
rect 11716 15484 11744 16374
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15638 11836 15982
rect 11992 15706 12020 16050
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11624 15456 11744 15484
rect 11980 15496 12032 15502
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 10966 14784 11022 14793
rect 10966 14719 11022 14728
rect 10980 13802 11008 14719
rect 11116 14716 11424 14736
rect 11116 14714 11122 14716
rect 11178 14714 11202 14716
rect 11258 14714 11282 14716
rect 11338 14714 11362 14716
rect 11418 14714 11424 14716
rect 11178 14662 11180 14714
rect 11360 14662 11362 14714
rect 11116 14660 11122 14662
rect 11178 14660 11202 14662
rect 11258 14660 11282 14662
rect 11338 14660 11362 14662
rect 11418 14660 11424 14662
rect 11116 14640 11424 14660
rect 11624 13802 11652 15456
rect 11980 15438 12032 15444
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11716 14006 11744 14282
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11808 13954 11836 14214
rect 11900 14074 11928 15302
rect 11992 14890 12020 15438
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14498 12020 14826
rect 12084 14618 12112 14962
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 11992 14482 12112 14498
rect 11992 14476 12124 14482
rect 11992 14470 12072 14476
rect 12072 14418 12124 14424
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11992 14006 12020 14350
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11980 14000 12032 14006
rect 11808 13926 11928 13954
rect 11980 13942 12032 13948
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 10980 12646 11008 13738
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11116 13628 11424 13648
rect 11116 13626 11122 13628
rect 11178 13626 11202 13628
rect 11258 13626 11282 13628
rect 11338 13626 11362 13628
rect 11418 13626 11424 13628
rect 11178 13574 11180 13626
rect 11360 13574 11362 13626
rect 11116 13572 11122 13574
rect 11178 13572 11202 13574
rect 11258 13572 11282 13574
rect 11338 13572 11362 13574
rect 11418 13572 11424 13574
rect 11116 13552 11424 13572
rect 11244 13320 11296 13326
rect 11296 13268 11468 13274
rect 11244 13262 11468 13268
rect 11256 13258 11468 13262
rect 11256 13252 11480 13258
rect 11256 13246 11428 13252
rect 11428 13194 11480 13200
rect 11716 12986 11744 13670
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11808 13394 11836 13466
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11116 12540 11424 12560
rect 11116 12538 11122 12540
rect 11178 12538 11202 12540
rect 11258 12538 11282 12540
rect 11338 12538 11362 12540
rect 11418 12538 11424 12540
rect 11178 12486 11180 12538
rect 11360 12486 11362 12538
rect 11116 12484 11122 12486
rect 11178 12484 11202 12486
rect 11258 12484 11282 12486
rect 11338 12484 11362 12486
rect 11418 12484 11424 12486
rect 11116 12464 11424 12484
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10506 9616 10562 9625
rect 10506 9551 10562 9560
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 9110 10456 9318
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10520 8974 10548 9551
rect 10612 9382 10640 10406
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 8968 10560 8974
rect 10428 8928 10508 8956
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10336 7886 10364 8842
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10428 7342 10456 8928
rect 10508 8910 10560 8916
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10416 7336 10468 7342
rect 10336 7296 10416 7324
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 7002 10180 7142
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10048 4684 10100 4690
rect 9784 4644 9904 4672
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9784 4078 9812 4490
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3738 9812 4014
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9678 3632 9734 3641
rect 9678 3567 9680 3576
rect 9732 3567 9734 3576
rect 9680 3538 9732 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 3058 9720 3334
rect 9784 3126 9812 3674
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9876 2990 9904 4644
rect 10048 4626 10100 4632
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3602 10088 4082
rect 10152 3738 10180 5510
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10060 3126 10088 3538
rect 10152 3398 10180 3674
rect 10244 3534 10272 7210
rect 10336 4146 10364 7296
rect 10416 7278 10468 7284
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 5710 10456 6802
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10520 4758 10548 7686
rect 10612 7410 10640 9318
rect 10704 9042 10732 10610
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10796 8974 10824 11086
rect 10888 10606 10916 11698
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11354 11008 11630
rect 11116 11452 11424 11472
rect 11116 11450 11122 11452
rect 11178 11450 11202 11452
rect 11258 11450 11282 11452
rect 11338 11450 11362 11452
rect 11418 11450 11424 11452
rect 11178 11398 11180 11450
rect 11360 11398 11362 11450
rect 11116 11396 11122 11398
rect 11178 11396 11202 11398
rect 11258 11396 11282 11398
rect 11338 11396 11362 11398
rect 11418 11396 11424 11398
rect 11116 11376 11424 11396
rect 11532 11354 11560 12582
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11624 11014 11652 12174
rect 11716 11898 11744 12271
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11116 10364 11424 10384
rect 11116 10362 11122 10364
rect 11178 10362 11202 10364
rect 11258 10362 11282 10364
rect 11338 10362 11362 10364
rect 11418 10362 11424 10364
rect 11178 10310 11180 10362
rect 11360 10310 11362 10362
rect 11116 10308 11122 10310
rect 11178 10308 11202 10310
rect 11258 10308 11282 10310
rect 11338 10308 11362 10310
rect 11418 10308 11424 10310
rect 11116 10288 11424 10308
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10888 9178 10916 9998
rect 11440 9586 11468 9998
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11116 9276 11424 9296
rect 11116 9274 11122 9276
rect 11178 9274 11202 9276
rect 11258 9274 11282 9276
rect 11338 9274 11362 9276
rect 11418 9274 11424 9276
rect 11178 9222 11180 9274
rect 11360 9222 11362 9274
rect 11116 9220 11122 9222
rect 11178 9220 11202 9222
rect 11258 9220 11282 9222
rect 11338 9220 11362 9222
rect 11418 9220 11424 9222
rect 11116 9200 11424 9220
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10888 8838 10916 9114
rect 11624 8974 11652 9930
rect 11716 9042 11744 10542
rect 11808 9450 11836 12854
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11612 8968 11664 8974
rect 10966 8936 11022 8945
rect 11612 8910 11664 8916
rect 10966 8871 11022 8880
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10980 8634 11008 8871
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 7546 10732 8366
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10796 7478 10824 8434
rect 11116 8188 11424 8208
rect 11116 8186 11122 8188
rect 11178 8186 11202 8188
rect 11258 8186 11282 8188
rect 11338 8186 11362 8188
rect 11418 8186 11424 8188
rect 11178 8134 11180 8186
rect 11360 8134 11362 8186
rect 11116 8132 11122 8134
rect 11178 8132 11202 8134
rect 11258 8132 11282 8134
rect 11338 8132 11362 8134
rect 11418 8132 11424 8134
rect 11116 8112 11424 8132
rect 11242 7984 11298 7993
rect 11242 7919 11298 7928
rect 11256 7886 11284 7919
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6390 10640 6598
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10704 6322 10732 6938
rect 10692 6316 10744 6322
rect 10796 6304 10824 7142
rect 10888 6458 10916 7822
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 7313 11192 7686
rect 11256 7410 11284 7822
rect 11244 7404 11296 7410
rect 11296 7364 11560 7392
rect 11244 7346 11296 7352
rect 11150 7304 11206 7313
rect 11150 7239 11206 7248
rect 11116 7100 11424 7120
rect 11116 7098 11122 7100
rect 11178 7098 11202 7100
rect 11258 7098 11282 7100
rect 11338 7098 11362 7100
rect 11418 7098 11424 7100
rect 11178 7046 11180 7098
rect 11360 7046 11362 7098
rect 11116 7044 11122 7046
rect 11178 7044 11202 7046
rect 11258 7044 11282 7046
rect 11338 7044 11362 7046
rect 11418 7044 11424 7046
rect 11116 7024 11424 7044
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10796 6276 10916 6304
rect 10692 6258 10744 6264
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10612 5778 10640 6122
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5166 10640 5714
rect 10704 5642 10732 6258
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10336 3126 10364 4082
rect 10428 3738 10456 4558
rect 10704 4554 10732 5578
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10796 4214 10824 6054
rect 10888 4282 10916 6276
rect 10980 6254 11008 6734
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5710 11008 6054
rect 11116 6012 11424 6032
rect 11116 6010 11122 6012
rect 11178 6010 11202 6012
rect 11258 6010 11282 6012
rect 11338 6010 11362 6012
rect 11418 6010 11424 6012
rect 11178 5958 11180 6010
rect 11360 5958 11362 6010
rect 11116 5956 11122 5958
rect 11178 5956 11202 5958
rect 11258 5956 11282 5958
rect 11338 5956 11362 5958
rect 11418 5956 11424 5958
rect 11116 5936 11424 5956
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11532 5234 11560 7364
rect 11624 6866 11652 8910
rect 11716 8294 11744 8978
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 7954 11744 8230
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11702 7848 11758 7857
rect 11702 7783 11704 7792
rect 11756 7783 11758 7792
rect 11704 7754 11756 7760
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11716 6798 11744 7754
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11624 6633 11652 6666
rect 11610 6624 11666 6633
rect 11610 6559 11666 6568
rect 11624 6322 11652 6559
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11624 5302 11652 6258
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11116 4924 11424 4944
rect 11116 4922 11122 4924
rect 11178 4922 11202 4924
rect 11258 4922 11282 4924
rect 11338 4922 11362 4924
rect 11418 4922 11424 4924
rect 11178 4870 11180 4922
rect 11360 4870 11362 4922
rect 11116 4868 11122 4870
rect 11178 4868 11202 4870
rect 11258 4868 11282 4870
rect 11338 4868 11362 4870
rect 11418 4868 11424 4870
rect 11116 4848 11424 4868
rect 11716 4622 11744 5646
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10520 3194 10548 3470
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 800 10180 2382
rect 10704 800 10732 3878
rect 11116 3836 11424 3856
rect 11116 3834 11122 3836
rect 11178 3834 11202 3836
rect 11258 3834 11282 3836
rect 11338 3834 11362 3836
rect 11418 3834 11424 3836
rect 11178 3782 11180 3834
rect 11360 3782 11362 3834
rect 11116 3780 11122 3782
rect 11178 3780 11202 3782
rect 11258 3780 11282 3782
rect 11338 3780 11362 3782
rect 11418 3780 11424 3782
rect 11116 3760 11424 3780
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10888 3126 10916 3402
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 11116 2748 11424 2768
rect 11116 2746 11122 2748
rect 11178 2746 11202 2748
rect 11258 2746 11282 2748
rect 11338 2746 11362 2748
rect 11418 2746 11424 2748
rect 11178 2694 11180 2746
rect 11360 2694 11362 2746
rect 11116 2692 11122 2694
rect 11178 2692 11202 2694
rect 11258 2692 11282 2694
rect 11338 2692 11362 2694
rect 11418 2692 11424 2694
rect 11116 2672 11424 2692
rect 11256 870 11376 898
rect 11256 800 11284 870
rect 7852 734 8156 762
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10690 0 10746 800
rect 11242 0 11298 800
rect 11348 762 11376 870
rect 11532 762 11560 3946
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3466 11652 3878
rect 11716 3738 11744 4014
rect 11808 3942 11836 8366
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11900 2774 11928 13926
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11992 12442 12020 13738
rect 12084 13734 12112 14282
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13326 12112 13670
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11762 12112 12174
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11980 9512 12032 9518
rect 11978 9480 11980 9489
rect 12032 9480 12034 9489
rect 11978 9415 12034 9424
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7410 12020 7890
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11992 6186 12020 6802
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11992 5710 12020 6122
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12084 5302 12112 11290
rect 12176 7002 12204 21830
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12360 21350 12388 21490
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12268 19174 12296 21286
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 20466 12480 20742
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12360 19553 12388 19654
rect 12346 19544 12402 19553
rect 12346 19479 12402 19488
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18630 12296 19110
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12360 17921 12388 18702
rect 12452 18272 12480 19178
rect 12544 18873 12572 20946
rect 12530 18864 12586 18873
rect 12530 18799 12586 18808
rect 12532 18284 12584 18290
rect 12452 18244 12532 18272
rect 12636 18272 12664 23990
rect 13004 23882 13032 23990
rect 13082 23911 13138 24711
rect 13634 23911 13690 24711
rect 14186 23911 14242 24711
rect 14738 23911 14794 24711
rect 15474 23911 15530 24711
rect 16026 23911 16082 24711
rect 16578 23911 16634 24711
rect 17130 23911 17186 24711
rect 17866 23911 17922 24711
rect 18418 23911 18474 24711
rect 18970 23911 19026 24711
rect 19522 23911 19578 24711
rect 20258 23911 20314 24711
rect 20810 23911 20866 24711
rect 21362 23911 21418 24711
rect 21914 23911 21970 24711
rect 22466 23911 22522 24711
rect 13096 23882 13124 23911
rect 13004 23854 13124 23882
rect 13648 22094 13676 23911
rect 13556 22066 13676 22094
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13268 21616 13320 21622
rect 13452 21616 13504 21622
rect 13320 21576 13452 21604
rect 13268 21558 13320 21564
rect 13452 21558 13504 21564
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 20466 12940 21286
rect 12900 20460 12952 20466
rect 12728 20420 12900 20448
rect 12728 19854 12756 20420
rect 12900 20402 12952 20408
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12898 20088 12954 20097
rect 12898 20023 12954 20032
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 19446 12756 19654
rect 12820 19446 12848 19477
rect 12716 19440 12768 19446
rect 12808 19440 12860 19446
rect 12716 19382 12768 19388
rect 12806 19408 12808 19417
rect 12860 19408 12862 19417
rect 12806 19343 12862 19352
rect 12636 18244 12756 18272
rect 12532 18226 12584 18232
rect 12346 17912 12402 17921
rect 12346 17847 12402 17856
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17542 12480 17682
rect 12544 17678 12572 18226
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 17882 12664 18090
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12346 17096 12402 17105
rect 12346 17031 12402 17040
rect 12360 16998 12388 17031
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 15638 12388 15982
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15162 12296 15302
rect 12452 15162 12480 16934
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12268 14278 12296 15098
rect 12544 15094 12572 15302
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12636 15026 12664 17818
rect 12728 17746 12756 18244
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12820 17105 12848 19343
rect 12912 18766 12940 20023
rect 13004 19242 13032 20402
rect 13096 19514 13124 21558
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 13188 21418 13216 21490
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 13280 20874 13308 21422
rect 13360 21140 13412 21146
rect 13464 21128 13492 21422
rect 13412 21100 13492 21128
rect 13360 21082 13412 21088
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13268 20868 13320 20874
rect 13268 20810 13320 20816
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13188 20330 13216 20810
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13188 19378 13216 20266
rect 13280 19854 13308 20402
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13372 19446 13400 20266
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 13004 18714 13032 19178
rect 13360 18896 13412 18902
rect 13174 18864 13230 18873
rect 13360 18838 13412 18844
rect 13230 18808 13308 18816
rect 13174 18799 13176 18808
rect 13228 18788 13308 18808
rect 13176 18770 13228 18776
rect 13004 18686 13124 18714
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12912 18290 12940 18566
rect 13004 18426 13032 18566
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 13096 18272 13124 18686
rect 13176 18284 13228 18290
rect 13096 18244 13176 18272
rect 13096 18086 13124 18244
rect 13176 18226 13228 18232
rect 13280 18170 13308 18788
rect 13188 18142 13308 18170
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13188 17134 13216 18142
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17338 13308 18022
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 17128 13228 17134
rect 12806 17096 12862 17105
rect 13176 17070 13228 17076
rect 12806 17031 12862 17040
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 15348 12756 16594
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15502 12848 16050
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15570 12940 15846
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12728 15320 12848 15348
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12268 13326 12296 13942
rect 12360 13802 12388 14894
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12360 13530 12388 13738
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12360 13025 12388 13194
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12452 12481 12480 14962
rect 12622 13424 12678 13433
rect 12820 13410 12848 15320
rect 12912 13938 12940 15370
rect 13004 14958 13032 16118
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12912 13530 12940 13874
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12820 13382 12940 13410
rect 12622 13359 12678 13368
rect 12636 13190 12664 13359
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12438 12472 12494 12481
rect 12438 12407 12440 12416
rect 12492 12407 12494 12416
rect 12440 12378 12492 12384
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12544 11801 12572 11834
rect 12254 11792 12310 11801
rect 12254 11727 12310 11736
rect 12530 11792 12586 11801
rect 12530 11727 12586 11736
rect 12268 11626 12296 11727
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 9586 12296 10950
rect 12360 10266 12388 11086
rect 12452 11082 12480 11494
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12636 10266 12664 12650
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12728 11354 12756 11698
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12820 10742 12848 12718
rect 12912 12306 12940 13382
rect 13188 12764 13216 17070
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13280 14414 13308 16186
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13268 12776 13320 12782
rect 13188 12736 13268 12764
rect 13268 12718 13320 12724
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11218 12940 11630
rect 13096 11558 13124 12106
rect 12992 11552 13044 11558
rect 12990 11520 12992 11529
rect 13084 11552 13136 11558
rect 13044 11520 13046 11529
rect 13084 11494 13136 11500
rect 12990 11455 13046 11464
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12360 9654 12388 10202
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12544 9586 12572 9998
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12268 9058 12296 9522
rect 12268 9042 12388 9058
rect 12256 9036 12388 9042
rect 12308 9030 12388 9036
rect 12256 8978 12308 8984
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7585 12296 7822
rect 12254 7576 12310 7585
rect 12254 7511 12256 7520
rect 12308 7511 12310 7520
rect 12256 7482 12308 7488
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6458 12204 6666
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4078 12112 4558
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12176 3738 12204 5510
rect 12268 4842 12296 7346
rect 12360 6633 12388 9030
rect 12544 8974 12572 9522
rect 12820 9489 12848 10678
rect 13004 10674 13032 11290
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 10198 13032 10610
rect 13082 10432 13138 10441
rect 13082 10367 13138 10376
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13004 10062 13032 10134
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13096 9926 13124 10367
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12806 9480 12862 9489
rect 12806 9415 12862 9424
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12452 8090 12480 8434
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12636 7886 12664 9318
rect 12728 8974 12756 9318
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12544 6798 12572 7754
rect 12636 7585 12664 7822
rect 12622 7576 12678 7585
rect 12622 7511 12678 7520
rect 12728 7410 12756 8910
rect 12820 8537 12848 9415
rect 12806 8528 12862 8537
rect 12806 8463 12862 8472
rect 12820 8430 12848 8463
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12820 7886 12848 7958
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12348 6384 12400 6390
rect 12452 6372 12480 6666
rect 12400 6344 12480 6372
rect 12348 6326 12400 6332
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12360 5098 12388 6054
rect 12544 5234 12572 6734
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 5778 12756 6598
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5370 12664 5510
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12912 5137 12940 7142
rect 12898 5128 12954 5137
rect 12348 5092 12400 5098
rect 12898 5063 12954 5072
rect 12348 5034 12400 5040
rect 12268 4814 12388 4842
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 3126 12020 3470
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11624 2746 11928 2774
rect 11624 2582 11652 2746
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12084 2514 12112 3538
rect 12176 3398 12204 3674
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 3040 12204 3334
rect 12268 3194 12296 4558
rect 12360 3602 12388 4814
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12636 4146 12664 4626
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12820 4146 12848 4490
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12636 3738 12664 4082
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12348 3596 12400 3602
rect 12400 3556 12572 3584
rect 12348 3538 12400 3544
rect 12438 3224 12494 3233
rect 12256 3188 12308 3194
rect 12544 3194 12572 3556
rect 12912 3534 12940 4150
rect 13004 3942 13032 4558
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 3233 12940 3470
rect 12898 3224 12954 3233
rect 12438 3159 12440 3168
rect 12256 3130 12308 3136
rect 12492 3159 12494 3168
rect 12532 3188 12584 3194
rect 12440 3130 12492 3136
rect 12898 3159 12954 3168
rect 12532 3130 12584 3136
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 12716 3052 12768 3058
rect 12176 3012 12716 3040
rect 12716 2994 12768 3000
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12440 2916 12492 2922
rect 12820 2904 12848 3062
rect 12492 2876 12848 2904
rect 12440 2858 12492 2864
rect 12176 2774 12204 2858
rect 12176 2746 12296 2774
rect 12268 2650 12296 2746
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11808 800 11836 2382
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12544 800 12572 2314
rect 13096 800 13124 3878
rect 13188 2310 13216 12582
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10266 13308 11086
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 7886 13308 8774
rect 13372 8514 13400 18838
rect 13464 17338 13492 20810
rect 13556 17377 13584 22066
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 21146 13676 21422
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13648 20806 13676 21082
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13740 20058 13768 21626
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 21010 13860 21490
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13726 19544 13782 19553
rect 13726 19479 13728 19488
rect 13780 19479 13782 19488
rect 13728 19450 13780 19456
rect 13832 19394 13860 20742
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13740 19366 13860 19394
rect 13740 17882 13768 19366
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13832 18290 13860 19246
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13542 17368 13598 17377
rect 13452 17332 13504 17338
rect 13542 17303 13598 17312
rect 13452 17274 13504 17280
rect 13648 16590 13676 17614
rect 13726 17096 13782 17105
rect 13726 17031 13782 17040
rect 13740 16726 13768 17031
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13832 16114 13860 17614
rect 13924 16522 13952 20402
rect 14016 19446 14044 20878
rect 14200 20534 14228 23911
rect 14752 22098 14780 23911
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14504 21788 14812 21808
rect 14504 21786 14510 21788
rect 14566 21786 14590 21788
rect 14646 21786 14670 21788
rect 14726 21786 14750 21788
rect 14806 21786 14812 21788
rect 14566 21734 14568 21786
rect 14748 21734 14750 21786
rect 14504 21732 14510 21734
rect 14566 21732 14590 21734
rect 14646 21732 14670 21734
rect 14726 21732 14750 21734
rect 14806 21732 14812 21734
rect 14504 21712 14812 21732
rect 14844 21690 14872 22170
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15108 22024 15160 22030
rect 14936 21984 15108 22012
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14370 21448 14426 21457
rect 14370 21383 14426 21392
rect 14384 21146 14412 21383
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14476 20874 14504 21558
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14504 20700 14812 20720
rect 14504 20698 14510 20700
rect 14566 20698 14590 20700
rect 14646 20698 14670 20700
rect 14726 20698 14750 20700
rect 14806 20698 14812 20700
rect 14566 20646 14568 20698
rect 14748 20646 14750 20698
rect 14504 20644 14510 20646
rect 14566 20644 14590 20646
rect 14646 20644 14670 20646
rect 14726 20644 14750 20646
rect 14806 20644 14812 20646
rect 14504 20624 14812 20644
rect 14844 20602 14872 20742
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14016 18766 14044 19382
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14016 17338 14044 17682
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16726 14044 17002
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15502 13676 15914
rect 14108 15910 14136 19722
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 19174 14228 19314
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14200 18154 14228 18906
rect 14384 18766 14412 20402
rect 14504 19612 14812 19632
rect 14504 19610 14510 19612
rect 14566 19610 14590 19612
rect 14646 19610 14670 19612
rect 14726 19610 14750 19612
rect 14806 19610 14812 19612
rect 14566 19558 14568 19610
rect 14748 19558 14750 19610
rect 14504 19556 14510 19558
rect 14566 19556 14590 19558
rect 14646 19556 14670 19558
rect 14726 19556 14750 19558
rect 14806 19556 14812 19558
rect 14504 19536 14812 19556
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14292 17882 14320 18566
rect 14384 18426 14412 18702
rect 14504 18524 14812 18544
rect 14504 18522 14510 18524
rect 14566 18522 14590 18524
rect 14646 18522 14670 18524
rect 14726 18522 14750 18524
rect 14806 18522 14812 18524
rect 14566 18470 14568 18522
rect 14748 18470 14750 18522
rect 14504 18468 14510 18470
rect 14566 18468 14590 18470
rect 14646 18468 14670 18470
rect 14726 18468 14750 18470
rect 14806 18468 14812 18470
rect 14504 18448 14812 18468
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14844 17882 14872 20402
rect 14936 19281 14964 21984
rect 15108 21966 15160 21972
rect 15396 21570 15424 22034
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15212 21542 15424 21570
rect 15028 21434 15056 21490
rect 15028 21406 15148 21434
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 20262 15056 21286
rect 15120 20942 15148 21406
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15120 20602 15148 20878
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 14922 19272 14978 19281
rect 14922 19207 14978 19216
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14936 18970 14964 19110
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14280 17876 14332 17882
rect 14200 17836 14280 17864
rect 14200 17202 14228 17836
rect 14280 17818 14332 17824
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14936 17746 14964 18566
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 15028 17678 15056 20198
rect 15120 18698 15148 20402
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15120 18290 15148 18634
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14504 17436 14812 17456
rect 14504 17434 14510 17436
rect 14566 17434 14590 17436
rect 14646 17434 14670 17436
rect 14726 17434 14750 17436
rect 14806 17434 14812 17436
rect 14566 17382 14568 17434
rect 14748 17382 14750 17434
rect 14504 17380 14510 17382
rect 14566 17380 14590 17382
rect 14646 17380 14670 17382
rect 14726 17380 14750 17382
rect 14806 17380 14812 17382
rect 14504 17360 14812 17380
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14186 16824 14242 16833
rect 14186 16759 14188 16768
rect 14240 16759 14242 16768
rect 14188 16730 14240 16736
rect 14292 16590 14320 17274
rect 14384 16794 14412 17274
rect 14844 16833 14872 17274
rect 14830 16824 14886 16833
rect 14372 16788 14424 16794
rect 14830 16759 14886 16768
rect 14372 16730 14424 16736
rect 15212 16674 15240 21542
rect 15488 21486 15516 23911
rect 16040 21622 16068 23911
rect 16592 22030 16620 23911
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15304 20466 15332 21422
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15304 17524 15332 20402
rect 15488 19854 15516 21286
rect 15856 21078 15884 21490
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 15844 21072 15896 21078
rect 15844 21014 15896 21020
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15488 19378 15516 19790
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18222 15516 18702
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 17678 15424 18022
rect 15474 17912 15530 17921
rect 15580 17882 15608 20810
rect 15856 20466 15884 21014
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15672 19718 15700 20334
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 20058 15792 20198
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15764 19514 15792 19994
rect 15856 19854 15884 20402
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15844 19372 15896 19378
rect 15764 19332 15844 19360
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 18766 15700 19110
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15672 18086 15700 18362
rect 15764 18222 15792 19332
rect 15844 19314 15896 19320
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15856 18766 15884 19178
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15660 18080 15712 18086
rect 15844 18080 15896 18086
rect 15660 18022 15712 18028
rect 15764 18040 15844 18068
rect 15474 17847 15530 17856
rect 15568 17876 15620 17882
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15304 17496 15424 17524
rect 15396 17202 15424 17496
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15304 16794 15332 17138
rect 15488 16998 15516 17847
rect 15568 17818 15620 17824
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15580 17202 15608 17546
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15476 16992 15528 16998
rect 15528 16952 15608 16980
rect 15476 16934 15528 16940
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 14372 16652 14424 16658
rect 15212 16646 15332 16674
rect 14372 16594 14424 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16182 14320 16526
rect 14384 16232 14412 16594
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14504 16348 14812 16368
rect 14504 16346 14510 16348
rect 14566 16346 14590 16348
rect 14646 16346 14670 16348
rect 14726 16346 14750 16348
rect 14806 16346 14812 16348
rect 14566 16294 14568 16346
rect 14748 16294 14750 16346
rect 14504 16292 14510 16294
rect 14566 16292 14590 16294
rect 14646 16292 14670 16294
rect 14726 16292 14750 16294
rect 14806 16292 14812 16294
rect 14504 16272 14812 16292
rect 14384 16204 14596 16232
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14568 16114 14596 16204
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14482 13492 14962
rect 13648 14822 13676 15438
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14074 13492 14418
rect 13648 14414 13676 14758
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13556 14278 13584 14350
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13464 11354 13492 12378
rect 13556 12238 13584 12650
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13556 10742 13584 12174
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13648 11150 13676 11562
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13556 9586 13584 10678
rect 13648 10606 13676 11086
rect 13832 10826 13860 15846
rect 14384 15502 14412 15846
rect 14568 15706 14596 16050
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14844 15570 14872 15846
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15026 14320 15302
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14016 14346 14044 14962
rect 14292 14618 14320 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14016 13938 14044 14282
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14016 13258 14044 13738
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14108 12986 14136 14554
rect 14384 14414 14412 15438
rect 14936 15434 14964 16458
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14504 15260 14812 15280
rect 14504 15258 14510 15260
rect 14566 15258 14590 15260
rect 14646 15258 14670 15260
rect 14726 15258 14750 15260
rect 14806 15258 14812 15260
rect 14566 15206 14568 15258
rect 14748 15206 14750 15258
rect 14504 15204 14510 15206
rect 14566 15204 14590 15206
rect 14646 15204 14670 15206
rect 14726 15204 14750 15206
rect 14806 15204 14812 15206
rect 14504 15184 14812 15204
rect 14936 15094 14964 15370
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14738 14512 14794 14521
rect 14738 14447 14740 14456
rect 14792 14447 14794 14456
rect 14740 14418 14792 14424
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14200 13530 14228 13942
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12850 14228 13466
rect 14292 13326 14320 14214
rect 14504 14172 14812 14192
rect 14504 14170 14510 14172
rect 14566 14170 14590 14172
rect 14646 14170 14670 14172
rect 14726 14170 14750 14172
rect 14806 14170 14812 14172
rect 14566 14118 14568 14170
rect 14748 14118 14750 14170
rect 14504 14116 14510 14118
rect 14566 14116 14590 14118
rect 14646 14116 14670 14118
rect 14726 14116 14750 14118
rect 14806 14116 14812 14118
rect 14504 14096 14812 14116
rect 14844 13938 14872 14214
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14936 13530 14964 15030
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12238 13952 12582
rect 14016 12442 14044 12786
rect 14384 12696 14412 13194
rect 14504 13084 14812 13104
rect 14504 13082 14510 13084
rect 14566 13082 14590 13084
rect 14646 13082 14670 13084
rect 14726 13082 14750 13084
rect 14806 13082 14812 13084
rect 14566 13030 14568 13082
rect 14748 13030 14750 13082
rect 14504 13028 14510 13030
rect 14566 13028 14590 13030
rect 14646 13028 14670 13030
rect 14726 13028 14750 13030
rect 14806 13028 14812 13030
rect 14504 13008 14812 13028
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14292 12668 14412 12696
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11218 14136 11494
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13832 10798 13952 10826
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13740 10266 13768 10474
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 10062 13860 10610
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13740 9518 13768 9862
rect 13832 9722 13860 9998
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13372 8486 13492 8514
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8090 13400 8230
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7970 13492 8486
rect 13372 7942 13492 7970
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 6390 13308 6734
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5710 13308 6190
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4146 13308 4966
rect 13372 4622 13400 7942
rect 13648 7546 13676 9454
rect 13740 8498 13768 9454
rect 13924 8634 13952 10798
rect 14200 10538 14228 12242
rect 14292 12238 14320 12668
rect 14752 12646 14780 12786
rect 14464 12640 14516 12646
rect 14462 12608 14464 12617
rect 14740 12640 14792 12646
rect 14516 12608 14518 12617
rect 14740 12582 14792 12588
rect 14462 12543 14518 12552
rect 14554 12472 14610 12481
rect 14554 12407 14610 12416
rect 14568 12306 14596 12407
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14752 12238 14780 12582
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14504 11996 14812 12016
rect 14504 11994 14510 11996
rect 14566 11994 14590 11996
rect 14646 11994 14670 11996
rect 14726 11994 14750 11996
rect 14806 11994 14812 11996
rect 14566 11942 14568 11994
rect 14748 11942 14750 11994
rect 14504 11940 14510 11942
rect 14566 11940 14590 11942
rect 14646 11940 14670 11942
rect 14726 11940 14750 11942
rect 14806 11940 14812 11942
rect 14504 11920 14812 11940
rect 14844 11762 14872 12174
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 11082 14596 11494
rect 14660 11286 14688 11698
rect 14830 11384 14886 11393
rect 14830 11319 14832 11328
rect 14884 11319 14886 11328
rect 14832 11290 14884 11296
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14504 10908 14812 10928
rect 14504 10906 14510 10908
rect 14566 10906 14590 10908
rect 14646 10906 14670 10908
rect 14726 10906 14750 10908
rect 14806 10906 14812 10908
rect 14566 10854 14568 10906
rect 14748 10854 14750 10906
rect 14504 10852 14510 10854
rect 14566 10852 14590 10854
rect 14646 10852 14670 10854
rect 14726 10852 14750 10854
rect 14806 10852 14812 10854
rect 14504 10832 14812 10852
rect 14844 10810 14872 11018
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 14016 9586 14044 9862
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13556 7274 13584 7346
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13464 6322 13492 6666
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13464 4146 13492 5102
rect 13556 5012 13584 7210
rect 13740 7206 13768 7686
rect 13924 7585 13952 7822
rect 13910 7576 13966 7585
rect 13910 7511 13966 7520
rect 13924 7410 13952 7511
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 6798 13768 7142
rect 13728 6792 13780 6798
rect 13648 6752 13728 6780
rect 13648 6322 13676 6752
rect 13728 6734 13780 6740
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5370 13676 5510
rect 13740 5370 13768 6054
rect 13832 5896 13860 7346
rect 14016 6118 14044 8570
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13832 5868 13952 5896
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13832 5166 13860 5714
rect 13924 5234 13952 5868
rect 14108 5710 14136 8774
rect 14200 8498 14228 10474
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 10266 14596 10406
rect 14556 10260 14608 10266
rect 14384 10220 14556 10248
rect 14384 9994 14412 10220
rect 14556 10202 14608 10208
rect 14660 9994 14688 10610
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14200 6186 14228 8434
rect 14292 6322 14320 9658
rect 14384 9654 14412 9930
rect 14504 9820 14812 9840
rect 14504 9818 14510 9820
rect 14566 9818 14590 9820
rect 14646 9818 14670 9820
rect 14726 9818 14750 9820
rect 14806 9818 14812 9820
rect 14566 9766 14568 9818
rect 14748 9766 14750 9818
rect 14504 9764 14510 9766
rect 14566 9764 14590 9766
rect 14646 9764 14670 9766
rect 14726 9764 14750 9766
rect 14806 9764 14812 9766
rect 14504 9744 14812 9764
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14384 8974 14412 9114
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14504 8732 14812 8752
rect 14504 8730 14510 8732
rect 14566 8730 14590 8732
rect 14646 8730 14670 8732
rect 14726 8730 14750 8732
rect 14806 8730 14812 8732
rect 14566 8678 14568 8730
rect 14748 8678 14750 8730
rect 14504 8676 14510 8678
rect 14566 8676 14590 8678
rect 14646 8676 14670 8678
rect 14726 8676 14750 8678
rect 14806 8676 14812 8678
rect 14504 8656 14812 8676
rect 14844 8566 14872 9318
rect 14936 8566 14964 13466
rect 15028 12986 15056 16118
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15106 13424 15162 13433
rect 15106 13359 15162 13368
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15028 12442 15056 12922
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15120 11830 15148 13359
rect 15212 12782 15240 13874
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15198 12608 15254 12617
rect 15198 12543 15254 12552
rect 15212 12442 15240 12543
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15304 11898 15332 16646
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15396 16250 15424 16526
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16250 15516 16390
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15580 16130 15608 16952
rect 15396 16102 15608 16130
rect 15396 12434 15424 16102
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15502 15608 15914
rect 15672 15910 15700 18022
rect 15764 16114 15792 18040
rect 15844 18022 15896 18028
rect 15948 17202 15976 19722
rect 16040 19378 16068 19994
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16132 18426 16160 20946
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16224 19334 16252 20470
rect 16408 20466 16436 21082
rect 16486 21040 16542 21049
rect 16486 20975 16542 20984
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19854 16344 20334
rect 16408 20058 16436 20402
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16500 19938 16528 20975
rect 16592 20602 16620 21354
rect 16762 21040 16818 21049
rect 16762 20975 16818 20984
rect 16776 20942 16804 20975
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16684 20466 16712 20742
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16408 19910 16528 19938
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19514 16344 19790
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16224 19306 16344 19334
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16040 18086 16068 18226
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 16040 17678 16068 17818
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15844 16992 15896 16998
rect 16040 16946 16068 17614
rect 15844 16934 15896 16940
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15764 16017 15792 16050
rect 15750 16008 15806 16017
rect 15750 15943 15806 15952
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14550 15516 14758
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15476 13320 15528 13326
rect 15474 13288 15476 13297
rect 15528 13288 15530 13297
rect 15474 13223 15530 13232
rect 15580 12594 15608 15098
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15672 13297 15700 14962
rect 15764 13938 15792 15943
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15750 13832 15806 13841
rect 15750 13767 15806 13776
rect 15658 13288 15714 13297
rect 15658 13223 15714 13232
rect 15580 12566 15700 12594
rect 15396 12406 15608 12434
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 15212 11014 15240 11834
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 11393 15332 11630
rect 15290 11384 15346 11393
rect 15396 11354 15424 11698
rect 15290 11319 15346 11328
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15292 11212 15344 11218
rect 15488 11200 15516 11290
rect 15344 11172 15516 11200
rect 15292 11154 15344 11160
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14370 8256 14426 8265
rect 14370 8191 14426 8200
rect 14384 6934 14412 8191
rect 14504 7644 14812 7664
rect 14504 7642 14510 7644
rect 14566 7642 14590 7644
rect 14646 7642 14670 7644
rect 14726 7642 14750 7644
rect 14806 7642 14812 7644
rect 14566 7590 14568 7642
rect 14748 7590 14750 7642
rect 14504 7588 14510 7590
rect 14566 7588 14590 7590
rect 14646 7588 14670 7590
rect 14726 7588 14750 7590
rect 14806 7588 14812 7590
rect 14504 7568 14812 7588
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14844 6730 14872 8298
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14936 7993 14964 8230
rect 14922 7984 14978 7993
rect 15028 7970 15056 9930
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 9178 15148 9522
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15120 8498 15148 8570
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15200 8424 15252 8430
rect 15106 8392 15162 8401
rect 15200 8366 15252 8372
rect 15106 8327 15108 8336
rect 15160 8327 15162 8336
rect 15108 8298 15160 8304
rect 15028 7942 15148 7970
rect 14922 7919 14978 7928
rect 14936 7410 14964 7919
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15028 6866 15056 7822
rect 15120 7342 15148 7942
rect 15212 7342 15240 8366
rect 15304 7886 15332 8774
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15120 6798 15148 7278
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13820 5160 13872 5166
rect 13818 5128 13820 5137
rect 13872 5128 13874 5137
rect 14200 5098 14228 6122
rect 14384 5778 14412 6598
rect 14504 6556 14812 6576
rect 14504 6554 14510 6556
rect 14566 6554 14590 6556
rect 14646 6554 14670 6556
rect 14726 6554 14750 6556
rect 14806 6554 14812 6556
rect 14566 6502 14568 6554
rect 14748 6502 14750 6554
rect 14504 6500 14510 6502
rect 14566 6500 14590 6502
rect 14646 6500 14670 6502
rect 14726 6500 14750 6502
rect 14806 6500 14812 6502
rect 14504 6480 14812 6500
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14384 5302 14412 5714
rect 14476 5710 14504 6122
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14660 5658 14688 6326
rect 14936 6322 14964 6598
rect 15028 6458 15056 6598
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15212 6202 15240 7278
rect 15396 7274 15424 9046
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 8090 15516 8434
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15488 7410 15516 7686
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 15120 6174 15240 6202
rect 14660 5630 14872 5658
rect 14504 5468 14812 5488
rect 14504 5466 14510 5468
rect 14566 5466 14590 5468
rect 14646 5466 14670 5468
rect 14726 5466 14750 5468
rect 14806 5466 14812 5468
rect 14566 5414 14568 5466
rect 14748 5414 14750 5466
rect 14504 5412 14510 5414
rect 14566 5412 14590 5414
rect 14646 5412 14670 5414
rect 14726 5412 14750 5414
rect 14806 5412 14812 5414
rect 14504 5392 14812 5412
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14738 5264 14794 5273
rect 14738 5199 14740 5208
rect 14792 5199 14794 5208
rect 14740 5170 14792 5176
rect 13818 5063 13874 5072
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 13636 5024 13688 5030
rect 13556 4984 13636 5012
rect 13636 4966 13688 4972
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13280 3670 13308 4082
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13280 3398 13308 3606
rect 13648 3534 13676 4966
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13648 3058 13676 3470
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13372 2514 13400 2994
rect 13832 2774 13860 4422
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 13912 3664 13964 3670
rect 13910 3632 13912 3641
rect 13964 3632 13966 3641
rect 13910 3567 13966 3576
rect 14292 3398 14320 3674
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14108 3194 14136 3334
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14384 3126 14412 4966
rect 14504 4380 14812 4400
rect 14504 4378 14510 4380
rect 14566 4378 14590 4380
rect 14646 4378 14670 4380
rect 14726 4378 14750 4380
rect 14806 4378 14812 4380
rect 14566 4326 14568 4378
rect 14748 4326 14750 4378
rect 14504 4324 14510 4326
rect 14566 4324 14590 4326
rect 14646 4324 14670 4326
rect 14726 4324 14750 4326
rect 14806 4324 14812 4326
rect 14504 4304 14812 4324
rect 14740 4072 14792 4078
rect 14844 4026 14872 5630
rect 14936 5234 14964 6122
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5778 15056 6054
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14792 4020 14872 4026
rect 14740 4014 14872 4020
rect 14752 3998 14872 4014
rect 14844 3534 14872 3998
rect 15028 3670 15056 5714
rect 15120 4146 15148 6174
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5030 15240 6054
rect 15304 5710 15332 7142
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4622 15240 4966
rect 15200 4616 15252 4622
rect 15252 4576 15332 4604
rect 15200 4558 15252 4564
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15212 4026 15240 4422
rect 15120 3998 15240 4026
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14504 3292 14812 3312
rect 14504 3290 14510 3292
rect 14566 3290 14590 3292
rect 14646 3290 14670 3292
rect 14726 3290 14750 3292
rect 14806 3290 14812 3292
rect 14566 3238 14568 3290
rect 14748 3238 14750 3290
rect 14504 3236 14510 3238
rect 14566 3236 14590 3238
rect 14646 3236 14670 3238
rect 14726 3236 14750 3238
rect 14806 3236 14812 3238
rect 14504 3216 14812 3236
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 15028 3058 15056 3606
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 13648 2746 13860 2774
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13372 2038 13400 2246
rect 13360 2032 13412 2038
rect 13360 1974 13412 1980
rect 13648 800 13676 2746
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14200 800 14228 2586
rect 15120 2258 15148 3998
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3534 15240 3878
rect 15304 3738 15332 4576
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15396 3534 15424 6695
rect 15488 6254 15516 7346
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 3534 15516 6190
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15396 3369 15424 3470
rect 15382 3360 15438 3369
rect 15382 3295 15438 3304
rect 15580 2582 15608 12406
rect 15672 12306 15700 12566
rect 15660 12300 15712 12306
rect 15764 12288 15792 13767
rect 15856 13258 15884 16934
rect 15948 16918 16068 16946
rect 15948 16590 15976 16918
rect 16132 16794 16160 17682
rect 16224 17678 16252 18294
rect 16316 17882 16344 19306
rect 16408 18086 16436 19910
rect 16488 19712 16540 19718
rect 16592 19700 16620 20198
rect 16540 19672 16620 19700
rect 16488 19654 16540 19660
rect 16500 19334 16528 19654
rect 16672 19372 16724 19378
rect 16500 19306 16620 19334
rect 16672 19314 16724 19320
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16408 17762 16436 18022
rect 16316 17734 16436 17762
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16120 16788 16172 16794
rect 16040 16748 16120 16776
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15948 12374 15976 16526
rect 16040 15162 16068 16748
rect 16120 16730 16172 16736
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16132 15026 16160 15438
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 16118 14920 16174 14929
rect 16040 14414 16068 14894
rect 16118 14855 16174 14864
rect 16132 14414 16160 14855
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16040 14074 16068 14350
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16132 13394 16160 14350
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16224 13274 16252 15846
rect 16040 13246 16252 13274
rect 16040 12442 16068 13246
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15764 12260 15884 12288
rect 15660 12242 15712 12248
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 11014 15700 11494
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 8945 15700 10610
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 8090 15700 8366
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15764 7750 15792 12106
rect 15856 11218 15884 12260
rect 16026 11520 16082 11529
rect 16026 11455 16082 11464
rect 16040 11286 16068 11455
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 8974 15884 10406
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8430 15884 8910
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15856 7886 15884 8366
rect 15948 8022 15976 10950
rect 16132 10742 16160 13126
rect 16224 12238 16252 13126
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16224 9994 16252 12174
rect 16316 11762 16344 17734
rect 16500 17610 16528 18702
rect 16592 18408 16620 19306
rect 16684 18902 16712 19314
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18970 16804 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16592 18380 16712 18408
rect 16578 18320 16634 18329
rect 16578 18255 16580 18264
rect 16632 18255 16634 18264
rect 16580 18226 16632 18232
rect 16580 17740 16632 17746
rect 16684 17728 16712 18380
rect 16776 18222 16804 18702
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17882 16804 18158
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16632 17700 16712 17728
rect 16580 17682 16632 17688
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16592 16697 16620 17138
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16578 16688 16634 16697
rect 16488 16652 16540 16658
rect 16578 16623 16634 16632
rect 16488 16594 16540 16600
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 15065 16436 16526
rect 16394 15056 16450 15065
rect 16394 14991 16450 15000
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16316 10810 16344 11086
rect 16408 11014 16436 14826
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16500 10826 16528 16594
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16114 16620 16390
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16684 15994 16712 17070
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16776 16590 16804 16730
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16592 15966 16712 15994
rect 16592 13394 16620 15966
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15570 16712 15846
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 15026 16712 15506
rect 16868 15042 16896 22034
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17052 21690 17080 21830
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16960 18970 16988 20946
rect 17144 20058 17172 23911
rect 17880 22506 17908 23911
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 17893 22332 18201 22352
rect 17893 22330 17899 22332
rect 17955 22330 17979 22332
rect 18035 22330 18059 22332
rect 18115 22330 18139 22332
rect 18195 22330 18201 22332
rect 17955 22278 17957 22330
rect 18137 22278 18139 22330
rect 17893 22276 17899 22278
rect 17955 22276 17979 22278
rect 18035 22276 18059 22278
rect 18115 22276 18139 22278
rect 18195 22276 18201 22278
rect 17893 22256 18201 22276
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17236 21350 17264 21830
rect 17420 21570 17448 22034
rect 17328 21542 17448 21570
rect 17500 21548 17552 21554
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17328 20618 17356 21542
rect 17500 21490 17552 21496
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17236 20590 17356 20618
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17236 19854 17264 20590
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 17224 19848 17276 19854
rect 17038 19816 17094 19825
rect 17224 19790 17276 19796
rect 17038 19751 17040 19760
rect 17092 19751 17094 19760
rect 17040 19722 17092 19728
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16960 18873 16988 18906
rect 16946 18864 17002 18873
rect 16946 18799 17002 18808
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16776 15014 16896 15042
rect 16776 14600 16804 15014
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 14618 16896 14894
rect 16684 14572 16804 14600
rect 16856 14612 16908 14618
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16408 10798 16528 10826
rect 16408 10441 16436 10798
rect 16488 10464 16540 10470
rect 16394 10432 16450 10441
rect 16488 10406 16540 10412
rect 16394 10367 16450 10376
rect 16500 10198 16528 10406
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 16040 7410 16068 8842
rect 16118 8528 16174 8537
rect 16118 8463 16120 8472
rect 16172 8463 16174 8472
rect 16120 8434 16172 8440
rect 16132 8022 16160 8434
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16028 7404 16080 7410
rect 15948 7364 16028 7392
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15752 7200 15804 7206
rect 15804 7160 15884 7188
rect 15752 7142 15804 7148
rect 15672 6934 15700 7142
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15660 6792 15712 6798
rect 15752 6792 15804 6798
rect 15660 6734 15712 6740
rect 15750 6760 15752 6769
rect 15804 6760 15806 6769
rect 15672 6633 15700 6734
rect 15750 6695 15806 6704
rect 15658 6624 15714 6633
rect 15658 6559 15714 6568
rect 15856 4146 15884 7160
rect 15948 4282 15976 7364
rect 16028 7346 16080 7352
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16040 6390 16068 6938
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 3534 15976 4082
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15672 3194 15700 3334
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 14936 2230 15148 2258
rect 14504 2204 14812 2224
rect 14504 2202 14510 2204
rect 14566 2202 14590 2204
rect 14646 2202 14670 2204
rect 14726 2202 14750 2204
rect 14806 2202 14812 2204
rect 14566 2150 14568 2202
rect 14748 2150 14750 2202
rect 14504 2148 14510 2150
rect 14566 2148 14590 2150
rect 14646 2148 14670 2150
rect 14726 2148 14750 2150
rect 14806 2148 14812 2150
rect 14504 2128 14812 2148
rect 14936 800 14964 2230
rect 15488 800 15516 2314
rect 16040 800 16068 5646
rect 16132 2990 16160 7958
rect 16316 7954 16344 9318
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16210 7304 16266 7313
rect 16210 7239 16266 7248
rect 16224 5302 16252 7239
rect 16316 7206 16344 7890
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 6118 16344 7142
rect 16408 6118 16436 8502
rect 16500 8498 16528 8910
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 7313 16528 7346
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16224 4826 16252 5102
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16316 2990 16344 5646
rect 16500 4690 16528 6938
rect 16592 6905 16620 12378
rect 16684 10996 16712 14572
rect 16856 14554 16908 14560
rect 16960 14498 16988 17614
rect 17052 16674 17080 18022
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17144 17134 17172 17682
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17236 16794 17264 19790
rect 17328 18290 17356 20470
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17314 16688 17370 16697
rect 17052 16646 17264 16674
rect 17040 16584 17092 16590
rect 17236 16561 17264 16646
rect 17314 16623 17370 16632
rect 17040 16526 17092 16532
rect 17222 16552 17278 16561
rect 17052 16046 17080 16526
rect 17222 16487 17278 16496
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 16182 17172 16390
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17052 15706 17080 15982
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14618 17172 14758
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16776 14470 16988 14498
rect 16776 11150 16804 14470
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16854 13968 16910 13977
rect 16854 13903 16910 13912
rect 16868 13394 16896 13903
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12594 16896 13126
rect 16960 12714 16988 14350
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 14074 17172 14214
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 12986 17080 13874
rect 17130 13424 17186 13433
rect 17130 13359 17186 13368
rect 17144 13326 17172 13359
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16868 12566 16988 12594
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16868 11898 16896 12174
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 11286 16896 11562
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16684 10968 16896 10996
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10169 16712 10610
rect 16670 10160 16726 10169
rect 16670 10095 16672 10104
rect 16724 10095 16726 10104
rect 16672 10066 16724 10072
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9110 16712 9930
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16684 8294 16712 9046
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16776 8090 16804 8978
rect 16868 8566 16896 10968
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16684 7818 16712 8026
rect 16776 7954 16804 8026
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16868 7410 16896 8502
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16868 6798 16896 7346
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5710 16620 6190
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16684 4706 16712 6258
rect 16776 5914 16804 6734
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16592 4678 16712 4706
rect 16592 4554 16620 4678
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 4282 16620 4490
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16684 4146 16712 4558
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3738 16620 4014
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16684 3670 16712 4082
rect 16776 3942 16804 5850
rect 16868 4622 16896 6598
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 4214 16896 4558
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16408 2854 16436 3402
rect 16868 2990 16896 4150
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16960 2774 16988 12566
rect 17052 9625 17080 12718
rect 17236 12646 17264 16487
rect 17328 14074 17356 16623
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17420 13682 17448 21354
rect 17512 20874 17540 21490
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17604 20942 17632 21354
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17788 21010 17816 21286
rect 17893 21244 18201 21264
rect 17893 21242 17899 21244
rect 17955 21242 17979 21244
rect 18035 21242 18059 21244
rect 18115 21242 18139 21244
rect 18195 21242 18201 21244
rect 17955 21190 17957 21242
rect 18137 21190 18139 21242
rect 17893 21188 17899 21190
rect 17955 21188 17979 21190
rect 18035 21188 18059 21190
rect 18115 21188 18139 21190
rect 18195 21188 18201 21190
rect 17893 21168 18201 21188
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17592 20936 17644 20942
rect 17880 20913 17908 20946
rect 17592 20878 17644 20884
rect 17866 20904 17922 20913
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 19446 17540 20810
rect 17604 20398 17632 20878
rect 17866 20839 17922 20848
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17696 20602 17724 20742
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17880 20244 17908 20839
rect 17696 20216 17908 20244
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17592 18828 17644 18834
rect 17696 18816 17724 20216
rect 17893 20156 18201 20176
rect 17893 20154 17899 20156
rect 17955 20154 17979 20156
rect 18035 20154 18059 20156
rect 18115 20154 18139 20156
rect 18195 20154 18201 20156
rect 17955 20102 17957 20154
rect 18137 20102 18139 20154
rect 17893 20100 17899 20102
rect 17955 20100 17979 20102
rect 18035 20100 18059 20102
rect 18115 20100 18139 20102
rect 18195 20100 18201 20102
rect 17893 20080 18201 20100
rect 18248 19922 18276 21490
rect 18340 19990 18368 22442
rect 18432 20058 18460 23911
rect 18694 23760 18750 23769
rect 18694 23695 18750 23704
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18524 22030 18552 22063
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 20942 18552 21286
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18524 20534 18552 20878
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 17788 18970 17816 19314
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 17893 19068 18201 19088
rect 17893 19066 17899 19068
rect 17955 19066 17979 19068
rect 18035 19066 18059 19068
rect 18115 19066 18139 19068
rect 18195 19066 18201 19068
rect 17955 19014 17957 19066
rect 18137 19014 18139 19066
rect 17893 19012 17899 19014
rect 17955 19012 17979 19014
rect 18035 19012 18059 19014
rect 18115 19012 18139 19014
rect 18195 19012 18201 19014
rect 17893 18992 18201 19012
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17644 18788 17724 18816
rect 17592 18770 17644 18776
rect 17498 17776 17554 17785
rect 17498 17711 17554 17720
rect 17512 17202 17540 17711
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16697 17540 17138
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 15162 17540 16526
rect 17604 16130 17632 18770
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 18426 17724 18566
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17788 18290 17816 18906
rect 18248 18766 18276 19110
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17893 17980 18201 18000
rect 17893 17978 17899 17980
rect 17955 17978 17979 17980
rect 18035 17978 18059 17980
rect 18115 17978 18139 17980
rect 18195 17978 18201 17980
rect 17955 17926 17957 17978
rect 18137 17926 18139 17978
rect 17893 17924 17899 17926
rect 17955 17924 17979 17926
rect 18035 17924 18059 17926
rect 18115 17924 18139 17926
rect 18195 17924 18201 17926
rect 17893 17904 18201 17924
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17682 17232 17738 17241
rect 17682 17167 17684 17176
rect 17736 17167 17738 17176
rect 17684 17138 17736 17144
rect 17696 16538 17724 17138
rect 17788 17105 17816 17478
rect 18156 17134 18184 17614
rect 18144 17128 18196 17134
rect 17774 17096 17830 17105
rect 18144 17070 18196 17076
rect 17774 17031 17830 17040
rect 17893 16892 18201 16912
rect 17893 16890 17899 16892
rect 17955 16890 17979 16892
rect 18035 16890 18059 16892
rect 18115 16890 18139 16892
rect 18195 16890 18201 16892
rect 17955 16838 17957 16890
rect 18137 16838 18139 16890
rect 17893 16836 17899 16838
rect 17955 16836 17979 16838
rect 18035 16836 18059 16838
rect 18115 16836 18139 16838
rect 18195 16836 18201 16838
rect 17893 16816 18201 16836
rect 18052 16720 18104 16726
rect 18248 16674 18276 18022
rect 18104 16668 18276 16674
rect 18052 16662 18276 16668
rect 18064 16646 18276 16662
rect 18064 16590 18092 16646
rect 18052 16584 18104 16590
rect 17696 16510 17816 16538
rect 18052 16526 18104 16532
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16250 17724 16390
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17604 16102 17724 16130
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15706 17632 15982
rect 17696 15978 17724 16102
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17512 14414 17540 14962
rect 17604 14822 17632 15370
rect 17696 15094 17724 15914
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17696 13938 17724 15030
rect 17788 14890 17816 16510
rect 17893 15804 18201 15824
rect 17893 15802 17899 15804
rect 17955 15802 17979 15804
rect 18035 15802 18059 15804
rect 18115 15802 18139 15804
rect 18195 15802 18201 15804
rect 17955 15750 17957 15802
rect 18137 15750 18139 15802
rect 17893 15748 17899 15750
rect 17955 15748 17979 15750
rect 18035 15748 18059 15750
rect 18115 15748 18139 15750
rect 18195 15748 18201 15750
rect 17893 15728 18201 15748
rect 18340 15502 18368 19246
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 17814 18460 18702
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18420 17672 18472 17678
rect 18524 17649 18552 19314
rect 18420 17614 18472 17620
rect 18510 17640 18566 17649
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17880 15026 17908 15438
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18248 15026 18276 15302
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17893 14716 18201 14736
rect 17893 14714 17899 14716
rect 17955 14714 17979 14716
rect 18035 14714 18059 14716
rect 18115 14714 18139 14716
rect 18195 14714 18201 14716
rect 17955 14662 17957 14714
rect 18137 14662 18139 14714
rect 17893 14660 17899 14662
rect 17955 14660 17979 14662
rect 18035 14660 18059 14662
rect 18115 14660 18139 14662
rect 18195 14660 18201 14662
rect 17893 14640 18201 14660
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 17420 13654 17632 13682
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17328 12442 17356 12786
rect 17420 12753 17448 12854
rect 17406 12744 17462 12753
rect 17406 12679 17462 12688
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17512 12322 17540 13466
rect 17328 12294 17540 12322
rect 17328 12238 17356 12294
rect 17316 12232 17368 12238
rect 17408 12232 17460 12238
rect 17316 12174 17368 12180
rect 17406 12200 17408 12209
rect 17460 12200 17462 12209
rect 17328 11608 17356 12174
rect 17406 12135 17462 12144
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17408 11620 17460 11626
rect 17328 11580 17408 11608
rect 17408 11562 17460 11568
rect 17314 11520 17370 11529
rect 17314 11455 17370 11464
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17038 9616 17094 9625
rect 17038 9551 17094 9560
rect 17144 9330 17172 11086
rect 17224 10464 17276 10470
rect 17222 10432 17224 10441
rect 17276 10432 17278 10441
rect 17222 10367 17278 10376
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17236 9450 17264 9930
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17144 9302 17264 9330
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17052 8362 17080 8910
rect 17144 8362 17172 8910
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 6866 17080 7822
rect 17144 7410 17172 8298
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17144 7313 17172 7346
rect 17130 7304 17186 7313
rect 17130 7239 17186 7248
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6769 17080 6802
rect 17038 6760 17094 6769
rect 17038 6695 17094 6704
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5370 17080 5510
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17144 3058 17172 6054
rect 17236 5914 17264 9302
rect 17328 6633 17356 11455
rect 17512 11150 17540 12038
rect 17604 11665 17632 13654
rect 17696 13258 17724 13738
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17788 12850 17816 14554
rect 18248 14414 18276 14962
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18142 13968 18198 13977
rect 18142 13903 18198 13912
rect 18156 13870 18184 13903
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18248 13734 18276 14010
rect 18340 13870 18368 14826
rect 18432 14464 18460 17614
rect 18510 17575 18566 17584
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16590 18552 17138
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18616 16114 18644 19722
rect 18708 18154 18736 23695
rect 18984 21962 19012 23911
rect 19246 22944 19302 22953
rect 19246 22879 19302 22888
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18800 18766 18828 20402
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18984 19310 19012 20198
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 19076 18442 19104 21490
rect 19154 21312 19210 21321
rect 19154 21247 19210 21256
rect 19168 19310 19196 21247
rect 19260 20602 19288 22879
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19352 19446 19380 21830
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19076 18414 19196 18442
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17134 18736 17614
rect 18800 17610 18828 18226
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18708 15706 18736 17070
rect 18800 17066 18828 17546
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18892 16998 18920 17138
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16046 18828 16526
rect 18892 16454 18920 16934
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18892 15502 18920 16390
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18432 14436 18644 14464
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 17893 13628 18201 13648
rect 17893 13626 17899 13628
rect 17955 13626 17979 13628
rect 18035 13626 18059 13628
rect 18115 13626 18139 13628
rect 18195 13626 18201 13628
rect 17955 13574 17957 13626
rect 18137 13574 18139 13626
rect 17893 13572 17899 13574
rect 17955 13572 17979 13574
rect 18035 13572 18059 13574
rect 18115 13572 18139 13574
rect 18195 13572 18201 13574
rect 17893 13552 18201 13572
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 13190 18092 13262
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17893 12540 18201 12560
rect 17893 12538 17899 12540
rect 17955 12538 17979 12540
rect 18035 12538 18059 12540
rect 18115 12538 18139 12540
rect 18195 12538 18201 12540
rect 17955 12486 17957 12538
rect 18137 12486 18139 12538
rect 17893 12484 17899 12486
rect 17955 12484 17979 12486
rect 18035 12484 18059 12486
rect 18115 12484 18139 12486
rect 18195 12484 18201 12486
rect 17893 12464 18201 12484
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17696 12345 17724 12378
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17696 11762 17724 12174
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17590 11656 17646 11665
rect 17590 11591 17646 11600
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11218 17632 11494
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17512 9722 17540 9930
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17314 6624 17370 6633
rect 17314 6559 17370 6568
rect 17328 6322 17356 6559
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17236 3602 17264 4762
rect 17420 4690 17448 9590
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17512 9489 17540 9522
rect 17498 9480 17554 9489
rect 17498 9415 17554 9424
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 9178 17540 9318
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8022 17540 8774
rect 17604 8514 17632 11018
rect 17696 10606 17724 11562
rect 17788 11354 17816 11698
rect 17880 11626 17908 12174
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11830 18184 12038
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18156 11694 18184 11766
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17893 11452 18201 11472
rect 17893 11450 17899 11452
rect 17955 11450 17979 11452
rect 18035 11450 18059 11452
rect 18115 11450 18139 11452
rect 18195 11450 18201 11452
rect 17955 11398 17957 11450
rect 18137 11398 18139 11450
rect 17893 11396 17899 11398
rect 17955 11396 17979 11398
rect 18035 11396 18059 11398
rect 18115 11396 18139 11398
rect 18195 11396 18201 11398
rect 17893 11376 18201 11396
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17788 10674 17816 11290
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17684 10600 17736 10606
rect 17736 10548 17816 10554
rect 17684 10542 17816 10548
rect 17696 10526 17816 10542
rect 17604 8486 17724 8514
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17512 7886 17540 7958
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17498 7576 17554 7585
rect 17498 7511 17554 7520
rect 17512 5166 17540 7511
rect 17604 5710 17632 8366
rect 17592 5704 17644 5710
rect 17696 5681 17724 8486
rect 17592 5646 17644 5652
rect 17682 5672 17738 5681
rect 17682 5607 17738 5616
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17500 5160 17552 5166
rect 17498 5128 17500 5137
rect 17552 5128 17554 5137
rect 17498 5063 17554 5072
rect 17592 5092 17644 5098
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4282 17448 4626
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17512 3398 17540 5063
rect 17592 5034 17644 5040
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17420 3126 17448 3334
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16960 2746 17172 2774
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16592 800 16620 2382
rect 16776 2038 16804 2586
rect 17144 2514 17172 2746
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16764 2032 16816 2038
rect 16764 1974 16816 1980
rect 11348 734 11560 762
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 16960 105 16988 2450
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 17328 800 17356 2314
rect 17604 921 17632 5034
rect 17696 4758 17724 5170
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17788 4604 17816 10526
rect 17893 10364 18201 10384
rect 17893 10362 17899 10364
rect 17955 10362 17979 10364
rect 18035 10362 18059 10364
rect 18115 10362 18139 10364
rect 18195 10362 18201 10364
rect 17955 10310 17957 10362
rect 18137 10310 18139 10362
rect 17893 10308 17899 10310
rect 17955 10308 17979 10310
rect 18035 10308 18059 10310
rect 18115 10308 18139 10310
rect 18195 10308 18201 10310
rect 17893 10288 18201 10308
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18248 10010 18276 13398
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18340 11762 18368 12786
rect 18432 12209 18460 14436
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18524 13734 18552 14282
rect 18616 14006 18644 14436
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18602 13288 18658 13297
rect 18512 13252 18564 13258
rect 18602 13223 18604 13232
rect 18512 13194 18564 13200
rect 18656 13223 18658 13232
rect 18604 13194 18656 13200
rect 18524 13161 18552 13194
rect 18510 13152 18566 13161
rect 18510 13087 18566 13096
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18418 12200 18474 12209
rect 18418 12135 18474 12144
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18524 10810 18552 11698
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18616 10742 18644 11698
rect 18708 11626 18736 12582
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 10736 18656 10742
rect 18708 10713 18736 11018
rect 18604 10678 18656 10684
rect 18694 10704 18750 10713
rect 18694 10639 18750 10648
rect 18064 9586 18092 9998
rect 18248 9982 18460 10010
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17893 9276 18201 9296
rect 17893 9274 17899 9276
rect 17955 9274 17979 9276
rect 18035 9274 18059 9276
rect 18115 9274 18139 9276
rect 18195 9274 18201 9276
rect 17955 9222 17957 9274
rect 18137 9222 18139 9274
rect 17893 9220 17899 9222
rect 17955 9220 17979 9222
rect 18035 9220 18059 9222
rect 18115 9220 18139 9222
rect 18195 9220 18201 9222
rect 17893 9200 18201 9220
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8634 18000 8774
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18156 8276 18184 8978
rect 18248 8974 18276 9862
rect 18326 9480 18382 9489
rect 18326 9415 18382 9424
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18340 8498 18368 9415
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18156 8248 18276 8276
rect 17893 8188 18201 8208
rect 17893 8186 17899 8188
rect 17955 8186 17979 8188
rect 18035 8186 18059 8188
rect 18115 8186 18139 8188
rect 18195 8186 18201 8188
rect 17955 8134 17957 8186
rect 18137 8134 18139 8186
rect 17893 8132 17899 8134
rect 17955 8132 17979 8134
rect 18035 8132 18059 8134
rect 18115 8132 18139 8134
rect 18195 8132 18201 8134
rect 17893 8112 18201 8132
rect 17958 7984 18014 7993
rect 17868 7948 17920 7954
rect 18248 7970 18276 8248
rect 17958 7919 18014 7928
rect 18156 7942 18276 7970
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 17868 7890 17920 7896
rect 17880 7546 17908 7890
rect 17972 7750 18000 7919
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 18156 7585 18184 7942
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18142 7576 18198 7585
rect 17868 7540 17920 7546
rect 18142 7511 18198 7520
rect 17868 7482 17920 7488
rect 18144 7404 18196 7410
rect 18248 7392 18276 7822
rect 18340 7546 18368 7958
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18196 7364 18276 7392
rect 18144 7346 18196 7352
rect 17893 7100 18201 7120
rect 17893 7098 17899 7100
rect 17955 7098 17979 7100
rect 18035 7098 18059 7100
rect 18115 7098 18139 7100
rect 18195 7098 18201 7100
rect 17955 7046 17957 7098
rect 18137 7046 18139 7098
rect 17893 7044 17899 7046
rect 17955 7044 17979 7046
rect 18035 7044 18059 7046
rect 18115 7044 18139 7046
rect 18195 7044 18201 7046
rect 17893 7024 18201 7044
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6322 18000 6598
rect 18248 6390 18276 7364
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 6769 18368 7346
rect 18432 7002 18460 9982
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18524 9178 18552 9522
rect 18616 9489 18644 9590
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18708 9110 18736 9590
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18708 8498 18736 9046
rect 18786 8528 18842 8537
rect 18696 8492 18748 8498
rect 18786 8463 18842 8472
rect 18696 8434 18748 8440
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 7886 18644 8298
rect 18800 7886 18828 8463
rect 18604 7880 18656 7886
rect 18788 7880 18840 7886
rect 18656 7840 18736 7868
rect 18604 7822 18656 7828
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18420 6792 18472 6798
rect 18326 6760 18382 6769
rect 18420 6734 18472 6740
rect 18326 6695 18382 6704
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17893 6012 18201 6032
rect 17893 6010 17899 6012
rect 17955 6010 17979 6012
rect 18035 6010 18059 6012
rect 18115 6010 18139 6012
rect 18195 6010 18201 6012
rect 17955 5958 17957 6010
rect 18137 5958 18139 6010
rect 17893 5956 17899 5958
rect 17955 5956 17979 5958
rect 18035 5956 18059 5958
rect 18115 5956 18139 5958
rect 18195 5956 18201 5958
rect 17893 5936 18201 5956
rect 18340 5166 18368 6598
rect 18432 6118 18460 6734
rect 18524 6322 18552 7686
rect 18616 7410 18644 7686
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 17893 4924 18201 4944
rect 17893 4922 17899 4924
rect 17955 4922 17979 4924
rect 18035 4922 18059 4924
rect 18115 4922 18139 4924
rect 18195 4922 18201 4924
rect 17955 4870 17957 4922
rect 18137 4870 18139 4922
rect 17893 4868 17899 4870
rect 17955 4868 17979 4870
rect 18035 4868 18059 4870
rect 18115 4868 18139 4870
rect 18195 4868 18201 4870
rect 17893 4848 18201 4868
rect 17696 4576 17816 4604
rect 17868 4616 17920 4622
rect 17696 2650 17724 4576
rect 17868 4558 17920 4564
rect 17880 4214 17908 4558
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 18248 4146 18276 4422
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17893 3836 18201 3856
rect 17893 3834 17899 3836
rect 17955 3834 17979 3836
rect 18035 3834 18059 3836
rect 18115 3834 18139 3836
rect 18195 3834 18201 3836
rect 17955 3782 17957 3834
rect 18137 3782 18139 3834
rect 17893 3780 17899 3782
rect 17955 3780 17979 3782
rect 18035 3780 18059 3782
rect 18115 3780 18139 3782
rect 18195 3780 18201 3782
rect 17893 3760 18201 3780
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17788 2530 17816 3674
rect 17958 3632 18014 3641
rect 17868 3596 17920 3602
rect 17958 3567 18014 3576
rect 17868 3538 17920 3544
rect 17880 3398 17908 3538
rect 17972 3534 18000 3567
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17868 3392 17920 3398
rect 18156 3369 18184 3470
rect 17868 3334 17920 3340
rect 18142 3360 18198 3369
rect 18142 3295 18198 3304
rect 18248 3194 18276 4082
rect 18432 3738 18460 5850
rect 18616 5778 18644 7142
rect 18708 6934 18736 7840
rect 18788 7822 18840 7828
rect 18800 7002 18828 7822
rect 18892 7562 18920 15438
rect 18984 12434 19012 18022
rect 19076 17785 19104 18226
rect 19062 17776 19118 17785
rect 19062 17711 19118 17720
rect 19168 16130 19196 18414
rect 19260 16697 19288 19314
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 17882 19380 18566
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19444 17762 19472 21422
rect 19536 20942 19564 23911
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19616 20800 19668 20806
rect 20180 20777 20208 21966
rect 19616 20742 19668 20748
rect 20166 20768 20222 20777
rect 19352 17734 19472 17762
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19352 17610 19380 17734
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17270 19472 17478
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19246 16688 19302 16697
rect 19246 16623 19302 16632
rect 19352 16590 19380 16934
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19168 16114 19288 16130
rect 19168 16108 19300 16114
rect 19168 16102 19248 16108
rect 19168 15502 19196 16102
rect 19248 16050 19300 16056
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19260 15881 19288 15914
rect 19246 15872 19302 15881
rect 19246 15807 19302 15816
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14249 19288 14826
rect 19352 14482 19380 15302
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19444 14618 19472 14962
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19246 14240 19302 14249
rect 19246 14175 19302 14184
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19260 13818 19288 13942
rect 19352 13938 19380 14418
rect 19536 13954 19564 17750
rect 19628 17626 19656 20742
rect 20166 20703 20222 20712
rect 20272 20534 20300 23911
rect 20628 20800 20680 20806
rect 20626 20768 20628 20777
rect 20680 20768 20682 20777
rect 20626 20703 20682 20712
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19720 19553 19748 20402
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19706 19544 19762 19553
rect 19706 19479 19762 19488
rect 19812 18970 19840 19722
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19417 19932 19654
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19812 18426 19840 18634
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 17678 20024 18226
rect 19984 17672 20036 17678
rect 19628 17598 19840 17626
rect 19984 17614 20036 17620
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19628 16794 19656 17478
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19720 16726 19748 17138
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19444 13926 19564 13954
rect 19260 13790 19380 13818
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18984 12406 19104 12434
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18984 11506 19012 11766
rect 19076 11608 19104 12406
rect 19168 11898 19196 12786
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19076 11580 19196 11608
rect 18984 11478 19104 11506
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18984 7750 19012 11086
rect 19076 10674 19104 11478
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19168 9674 19196 11580
rect 19260 11529 19288 12038
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19352 11218 19380 13790
rect 19444 13734 19472 13926
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19536 13326 19564 13738
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12986 19472 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19536 11898 19564 12310
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10742 19380 10950
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19352 10062 19380 10678
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19076 9646 19196 9674
rect 19076 8401 19104 9646
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 8537 19196 8570
rect 19154 8528 19210 8537
rect 19154 8463 19156 8472
rect 19208 8463 19210 8472
rect 19156 8434 19208 8440
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18892 7534 19012 7562
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18708 6798 18736 6870
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18786 6760 18842 6769
rect 18786 6695 18842 6704
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18708 5914 18736 6190
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18524 5098 18552 5646
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18524 4826 18552 5034
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18616 4690 18644 5714
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18708 5370 18736 5578
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18708 4622 18736 5306
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 3058 18276 3130
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 17893 2748 18201 2768
rect 17893 2746 17899 2748
rect 17955 2746 17979 2748
rect 18035 2746 18059 2748
rect 18115 2746 18139 2748
rect 18195 2746 18201 2748
rect 17955 2694 17957 2746
rect 18137 2694 18139 2746
rect 17893 2692 17899 2694
rect 17955 2692 17979 2694
rect 18035 2692 18059 2694
rect 18115 2692 18139 2694
rect 18195 2692 18201 2694
rect 17893 2672 18201 2692
rect 17788 2502 17908 2530
rect 17590 912 17646 921
rect 17590 847 17646 856
rect 17880 800 17908 2502
rect 18340 1714 18368 3334
rect 18432 2990 18460 3674
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18616 2514 18644 3606
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18800 2310 18828 6695
rect 18892 6225 18920 7346
rect 18878 6216 18934 6225
rect 18878 6151 18934 6160
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 2553 18920 5510
rect 18878 2544 18934 2553
rect 18984 2530 19012 7534
rect 19076 7478 19104 7822
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19168 7410 19196 8230
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19168 6934 19196 7346
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 5302 19104 6734
rect 19168 6730 19196 6870
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 19260 6168 19288 9454
rect 19444 8090 19472 11086
rect 19536 10606 19564 11494
rect 19628 10674 19656 14350
rect 19720 14006 19748 15030
rect 19812 14074 19840 17598
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19904 15065 19932 15438
rect 19890 15056 19946 15065
rect 19890 14991 19946 15000
rect 19996 14074 20024 17614
rect 20088 17338 20116 20198
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20456 18601 20484 19790
rect 20628 19712 20680 19718
rect 20626 19680 20628 19689
rect 20680 19680 20682 19689
rect 20626 19615 20682 19624
rect 20824 19242 20852 23911
rect 21376 22098 21404 23911
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21928 20942 21956 23911
rect 22480 21554 22508 23911
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20640 18714 20668 18770
rect 20640 18686 20760 18714
rect 20442 18592 20498 18601
rect 20442 18527 20498 18536
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20272 18086 20300 18362
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20272 17338 20300 18022
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20456 17202 20484 17750
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20548 17202 20576 17614
rect 20640 17338 20668 17614
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 17218 20760 18686
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20640 17190 20760 17218
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 15162 20116 16934
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20088 14414 20116 15098
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19720 12238 19748 13466
rect 19812 12442 19840 13670
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19904 12170 19932 13874
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19996 12646 20024 12922
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12442 20024 12582
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19536 10266 19564 10542
rect 19628 10470 19656 10610
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19812 9602 19840 11154
rect 20088 11098 20116 14350
rect 20180 13938 20208 15438
rect 20272 14346 20300 15982
rect 20364 15094 20392 16594
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20456 15162 20484 15846
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20180 11830 20208 12854
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20272 11694 20300 14282
rect 20456 14074 20484 14758
rect 20548 14414 20576 16050
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20364 12850 20392 13806
rect 20456 13462 20484 14010
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 13530 20576 13874
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20456 12730 20484 13398
rect 20640 13394 20668 17190
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20732 14618 20760 15914
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20364 12702 20484 12730
rect 20364 12238 20392 12702
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12306 20668 12582
rect 20732 12345 20760 13194
rect 20718 12336 20774 12345
rect 20628 12300 20680 12306
rect 20718 12271 20774 12280
rect 20628 12242 20680 12248
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19904 11070 20116 11098
rect 19904 10470 19932 11070
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19996 10810 20024 10950
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10266 19932 10406
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19996 10198 20024 10542
rect 20088 10266 20116 10950
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 20272 10130 20300 11630
rect 20548 10674 20576 11766
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20640 10606 20668 12242
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20640 10062 20668 10406
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 19812 9574 19932 9602
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 8974 19748 9318
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19812 8838 19840 9386
rect 19904 9042 19932 9574
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19800 8832 19852 8838
rect 20732 8809 20760 8842
rect 19800 8774 19852 8780
rect 20718 8800 20774 8809
rect 19536 8498 19564 8774
rect 20718 8735 20774 8744
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 6866 19380 7686
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19168 6140 19288 6168
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19168 5166 19196 6140
rect 19246 6080 19302 6089
rect 19246 6015 19302 6024
rect 19260 5914 19288 6015
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19338 5808 19394 5817
rect 19338 5743 19394 5752
rect 19352 5710 19380 5743
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19444 5302 19472 6598
rect 19536 6322 19564 7958
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19168 4282 19196 4422
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19168 4146 19196 4218
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19168 2650 19196 4082
rect 19352 4078 19380 4558
rect 19444 4554 19472 5238
rect 19812 4826 19840 6394
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 19628 4214 19656 4490
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3602 19380 4014
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19720 3534 19748 4082
rect 19708 3528 19760 3534
rect 19522 3496 19578 3505
rect 19708 3470 19760 3476
rect 19522 3431 19524 3440
rect 19576 3431 19578 3440
rect 19524 3402 19576 3408
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 18984 2502 19104 2530
rect 18878 2479 18934 2488
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18340 1686 18460 1714
rect 18432 800 18460 1686
rect 18984 800 19012 2382
rect 19076 2106 19104 2502
rect 19064 2100 19116 2106
rect 19064 2042 19116 2048
rect 19720 800 19748 2994
rect 19904 2038 19932 7142
rect 20180 7002 20208 7278
rect 20272 7274 20300 8026
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20088 6118 20116 6734
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19982 5944 20038 5953
rect 19982 5879 19984 5888
rect 20036 5879 20038 5888
rect 19984 5850 20036 5856
rect 20088 3942 20116 6054
rect 20180 5574 20208 6122
rect 20272 5778 20300 7210
rect 20548 7177 20576 7754
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20534 7168 20590 7177
rect 20534 7103 20590 7112
rect 20640 6662 20668 7686
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20364 5370 20392 5646
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20548 5273 20576 6258
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5846 20668 6054
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20534 5264 20590 5273
rect 20534 5199 20590 5208
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20732 4457 20760 4490
rect 20718 4448 20774 4457
rect 20718 4383 20774 4392
rect 20258 4176 20314 4185
rect 20258 4111 20260 4120
rect 20312 4111 20314 4120
rect 20260 4082 20312 4088
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19892 2032 19944 2038
rect 19892 1974 19944 1980
rect 19996 1737 20024 3402
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 19982 1728 20038 1737
rect 19982 1663 20038 1672
rect 20272 800 20300 2994
rect 20824 800 20852 3946
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 800 21404 3878
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21928 800 21956 3402
rect 16946 96 17002 105
rect 16946 31 17002 40
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
<< via2 >>
rect 3146 24520 3202 24576
rect 1582 20168 1638 20224
rect 1858 22072 1914 22128
rect 1398 19352 1454 19408
rect 1674 18536 1730 18592
rect 2318 22888 2374 22944
rect 2318 19372 2374 19408
rect 2318 19352 2320 19372
rect 2320 19352 2372 19372
rect 2372 19352 2374 19372
rect 1858 17448 1914 17504
rect 1398 15000 1454 15056
rect 1674 13912 1730 13968
rect 1582 13096 1638 13152
rect 1214 10104 1270 10160
rect 1582 11500 1584 11520
rect 1584 11500 1636 11520
rect 1636 11500 1638 11520
rect 1582 11464 1638 11500
rect 1582 10412 1584 10432
rect 1584 10412 1636 10432
rect 1636 10412 1638 10432
rect 1582 10376 1638 10412
rect 1858 12280 1914 12336
rect 2778 23704 2834 23760
rect 4344 22330 4400 22332
rect 4424 22330 4480 22332
rect 4504 22330 4560 22332
rect 4584 22330 4640 22332
rect 4344 22278 4390 22330
rect 4390 22278 4400 22330
rect 4424 22278 4454 22330
rect 4454 22278 4466 22330
rect 4466 22278 4480 22330
rect 4504 22278 4518 22330
rect 4518 22278 4530 22330
rect 4530 22278 4560 22330
rect 4584 22278 4594 22330
rect 4594 22278 4640 22330
rect 4344 22276 4400 22278
rect 4424 22276 4480 22278
rect 4504 22276 4560 22278
rect 4584 22276 4640 22278
rect 3238 20984 3294 21040
rect 3330 17176 3386 17232
rect 2686 15952 2742 16008
rect 2778 15816 2834 15872
rect 1766 9560 1822 9616
rect 1674 8336 1730 8392
rect 1674 7928 1730 7984
rect 1950 8780 1952 8800
rect 1952 8780 2004 8800
rect 2004 8780 2006 8800
rect 1950 8744 2006 8780
rect 2778 15000 2834 15056
rect 3514 15000 3570 15056
rect 1858 6840 1914 6896
rect 2226 6840 2282 6896
rect 1766 6568 1822 6624
rect 1950 6024 2006 6080
rect 1858 5652 1860 5672
rect 1860 5652 1912 5672
rect 1912 5652 1914 5672
rect 1858 5616 1914 5652
rect 2042 5228 2098 5264
rect 2042 5208 2044 5228
rect 2044 5208 2096 5228
rect 2096 5208 2098 5228
rect 1398 4392 1454 4448
rect 1858 856 1914 912
rect 2778 2488 2834 2544
rect 4344 21242 4400 21244
rect 4424 21242 4480 21244
rect 4504 21242 4560 21244
rect 4584 21242 4640 21244
rect 4344 21190 4390 21242
rect 4390 21190 4400 21242
rect 4424 21190 4454 21242
rect 4454 21190 4466 21242
rect 4466 21190 4480 21242
rect 4504 21190 4518 21242
rect 4518 21190 4530 21242
rect 4530 21190 4560 21242
rect 4584 21190 4594 21242
rect 4594 21190 4640 21242
rect 4344 21188 4400 21190
rect 4424 21188 4480 21190
rect 4504 21188 4560 21190
rect 4584 21188 4640 21190
rect 4344 20154 4400 20156
rect 4424 20154 4480 20156
rect 4504 20154 4560 20156
rect 4584 20154 4640 20156
rect 4344 20102 4390 20154
rect 4390 20102 4400 20154
rect 4424 20102 4454 20154
rect 4454 20102 4466 20154
rect 4466 20102 4480 20154
rect 4504 20102 4518 20154
rect 4518 20102 4530 20154
rect 4530 20102 4560 20154
rect 4584 20102 4594 20154
rect 4594 20102 4640 20154
rect 4344 20100 4400 20102
rect 4424 20100 4480 20102
rect 4504 20100 4560 20102
rect 4584 20100 4640 20102
rect 3882 19236 3938 19272
rect 3882 19216 3884 19236
rect 3884 19216 3936 19236
rect 3936 19216 3938 19236
rect 4250 19216 4306 19272
rect 4344 19066 4400 19068
rect 4424 19066 4480 19068
rect 4504 19066 4560 19068
rect 4584 19066 4640 19068
rect 4344 19014 4390 19066
rect 4390 19014 4400 19066
rect 4424 19014 4454 19066
rect 4454 19014 4466 19066
rect 4466 19014 4480 19066
rect 4504 19014 4518 19066
rect 4518 19014 4530 19066
rect 4530 19014 4560 19066
rect 4584 19014 4594 19066
rect 4594 19014 4640 19066
rect 4344 19012 4400 19014
rect 4424 19012 4480 19014
rect 4504 19012 4560 19014
rect 4584 19012 4640 19014
rect 4066 17584 4122 17640
rect 4344 17978 4400 17980
rect 4424 17978 4480 17980
rect 4504 17978 4560 17980
rect 4584 17978 4640 17980
rect 4344 17926 4390 17978
rect 4390 17926 4400 17978
rect 4424 17926 4454 17978
rect 4454 17926 4466 17978
rect 4466 17926 4480 17978
rect 4504 17926 4518 17978
rect 4518 17926 4530 17978
rect 4530 17926 4560 17978
rect 4584 17926 4594 17978
rect 4594 17926 4640 17978
rect 4344 17924 4400 17926
rect 4424 17924 4480 17926
rect 4504 17924 4560 17926
rect 4584 17924 4640 17926
rect 4344 16890 4400 16892
rect 4424 16890 4480 16892
rect 4504 16890 4560 16892
rect 4584 16890 4640 16892
rect 4344 16838 4390 16890
rect 4390 16838 4400 16890
rect 4424 16838 4454 16890
rect 4454 16838 4466 16890
rect 4466 16838 4480 16890
rect 4504 16838 4518 16890
rect 4518 16838 4530 16890
rect 4530 16838 4560 16890
rect 4584 16838 4594 16890
rect 4594 16838 4640 16890
rect 4344 16836 4400 16838
rect 4424 16836 4480 16838
rect 4504 16836 4560 16838
rect 4584 16836 4640 16838
rect 4066 16632 4122 16688
rect 4802 19352 4858 19408
rect 5354 20440 5410 20496
rect 5354 20340 5356 20360
rect 5356 20340 5408 20360
rect 5408 20340 5410 20360
rect 5354 20304 5410 20340
rect 5814 20576 5870 20632
rect 4344 15802 4400 15804
rect 4424 15802 4480 15804
rect 4504 15802 4560 15804
rect 4584 15802 4640 15804
rect 4344 15750 4390 15802
rect 4390 15750 4400 15802
rect 4424 15750 4454 15802
rect 4454 15750 4466 15802
rect 4466 15750 4480 15802
rect 4504 15750 4518 15802
rect 4518 15750 4530 15802
rect 4530 15750 4560 15802
rect 4584 15750 4594 15802
rect 4594 15750 4640 15802
rect 4344 15748 4400 15750
rect 4424 15748 4480 15750
rect 4504 15748 4560 15750
rect 4584 15748 4640 15750
rect 4344 14714 4400 14716
rect 4424 14714 4480 14716
rect 4504 14714 4560 14716
rect 4584 14714 4640 14716
rect 4344 14662 4390 14714
rect 4390 14662 4400 14714
rect 4424 14662 4454 14714
rect 4454 14662 4466 14714
rect 4466 14662 4480 14714
rect 4504 14662 4518 14714
rect 4518 14662 4530 14714
rect 4530 14662 4560 14714
rect 4584 14662 4594 14714
rect 4594 14662 4640 14714
rect 4344 14660 4400 14662
rect 4424 14660 4480 14662
rect 4504 14660 4560 14662
rect 4584 14660 4640 14662
rect 4344 13626 4400 13628
rect 4424 13626 4480 13628
rect 4504 13626 4560 13628
rect 4584 13626 4640 13628
rect 4344 13574 4390 13626
rect 4390 13574 4400 13626
rect 4424 13574 4454 13626
rect 4454 13574 4466 13626
rect 4466 13574 4480 13626
rect 4504 13574 4518 13626
rect 4518 13574 4530 13626
rect 4530 13574 4560 13626
rect 4584 13574 4594 13626
rect 4594 13574 4640 13626
rect 4344 13572 4400 13574
rect 4424 13572 4480 13574
rect 4504 13572 4560 13574
rect 4584 13572 4640 13574
rect 4344 12538 4400 12540
rect 4424 12538 4480 12540
rect 4504 12538 4560 12540
rect 4584 12538 4640 12540
rect 4344 12486 4390 12538
rect 4390 12486 4400 12538
rect 4424 12486 4454 12538
rect 4454 12486 4466 12538
rect 4466 12486 4480 12538
rect 4504 12486 4518 12538
rect 4518 12486 4530 12538
rect 4530 12486 4560 12538
rect 4584 12486 4594 12538
rect 4594 12486 4640 12538
rect 4344 12484 4400 12486
rect 4424 12484 4480 12486
rect 4504 12484 4560 12486
rect 4584 12484 4640 12486
rect 3974 12280 4030 12336
rect 4344 11450 4400 11452
rect 4424 11450 4480 11452
rect 4504 11450 4560 11452
rect 4584 11450 4640 11452
rect 4344 11398 4390 11450
rect 4390 11398 4400 11450
rect 4424 11398 4454 11450
rect 4454 11398 4466 11450
rect 4466 11398 4480 11450
rect 4504 11398 4518 11450
rect 4518 11398 4530 11450
rect 4530 11398 4560 11450
rect 4584 11398 4594 11450
rect 4594 11398 4640 11450
rect 4344 11396 4400 11398
rect 4424 11396 4480 11398
rect 4504 11396 4560 11398
rect 4584 11396 4640 11398
rect 6090 20304 6146 20360
rect 6274 20476 6276 20496
rect 6276 20476 6328 20496
rect 6328 20476 6330 20496
rect 6274 20440 6330 20476
rect 5722 14764 5724 14784
rect 5724 14764 5776 14784
rect 5776 14764 5778 14784
rect 5722 14728 5778 14764
rect 5814 14048 5870 14104
rect 4344 10362 4400 10364
rect 4424 10362 4480 10364
rect 4504 10362 4560 10364
rect 4584 10362 4640 10364
rect 4344 10310 4390 10362
rect 4390 10310 4400 10362
rect 4424 10310 4454 10362
rect 4454 10310 4466 10362
rect 4466 10310 4480 10362
rect 4504 10310 4518 10362
rect 4518 10310 4530 10362
rect 4530 10310 4560 10362
rect 4584 10310 4594 10362
rect 4594 10310 4640 10362
rect 4344 10308 4400 10310
rect 4424 10308 4480 10310
rect 4504 10308 4560 10310
rect 4584 10308 4640 10310
rect 4344 9274 4400 9276
rect 4424 9274 4480 9276
rect 4504 9274 4560 9276
rect 4584 9274 4640 9276
rect 4344 9222 4390 9274
rect 4390 9222 4400 9274
rect 4424 9222 4454 9274
rect 4454 9222 4466 9274
rect 4466 9222 4480 9274
rect 4504 9222 4518 9274
rect 4518 9222 4530 9274
rect 4530 9222 4560 9274
rect 4584 9222 4594 9274
rect 4594 9222 4640 9274
rect 4344 9220 4400 9222
rect 4424 9220 4480 9222
rect 4504 9220 4560 9222
rect 4584 9220 4640 9222
rect 4158 9016 4214 9072
rect 3514 7928 3570 7984
rect 3698 7792 3754 7848
rect 4344 8186 4400 8188
rect 4424 8186 4480 8188
rect 4504 8186 4560 8188
rect 4584 8186 4640 8188
rect 4344 8134 4390 8186
rect 4390 8134 4400 8186
rect 4424 8134 4454 8186
rect 4454 8134 4466 8186
rect 4466 8134 4480 8186
rect 4504 8134 4518 8186
rect 4518 8134 4530 8186
rect 4530 8134 4560 8186
rect 4584 8134 4594 8186
rect 4594 8134 4640 8186
rect 4344 8132 4400 8134
rect 4424 8132 4480 8134
rect 4504 8132 4560 8134
rect 4584 8132 4640 8134
rect 4344 7098 4400 7100
rect 4424 7098 4480 7100
rect 4504 7098 4560 7100
rect 4584 7098 4640 7100
rect 4344 7046 4390 7098
rect 4390 7046 4400 7098
rect 4424 7046 4454 7098
rect 4454 7046 4466 7098
rect 4466 7046 4480 7098
rect 4504 7046 4518 7098
rect 4518 7046 4530 7098
rect 4530 7046 4560 7098
rect 4584 7046 4594 7098
rect 4594 7046 4640 7098
rect 4344 7044 4400 7046
rect 4424 7044 4480 7046
rect 4504 7044 4560 7046
rect 4584 7044 4640 7046
rect 4344 6010 4400 6012
rect 4424 6010 4480 6012
rect 4504 6010 4560 6012
rect 4584 6010 4640 6012
rect 4344 5958 4390 6010
rect 4390 5958 4400 6010
rect 4424 5958 4454 6010
rect 4454 5958 4466 6010
rect 4466 5958 4480 6010
rect 4504 5958 4518 6010
rect 4518 5958 4530 6010
rect 4530 5958 4560 6010
rect 4584 5958 4594 6010
rect 4594 5958 4640 6010
rect 4344 5956 4400 5958
rect 4424 5956 4480 5958
rect 4504 5956 4560 5958
rect 4584 5956 4640 5958
rect 4344 4922 4400 4924
rect 4424 4922 4480 4924
rect 4504 4922 4560 4924
rect 4584 4922 4640 4924
rect 4344 4870 4390 4922
rect 4390 4870 4400 4922
rect 4424 4870 4454 4922
rect 4454 4870 4466 4922
rect 4466 4870 4480 4922
rect 4504 4870 4518 4922
rect 4518 4870 4530 4922
rect 4530 4870 4560 4922
rect 4584 4870 4594 4922
rect 4594 4870 4640 4922
rect 4344 4868 4400 4870
rect 4424 4868 4480 4870
rect 4504 4868 4560 4870
rect 4584 4868 4640 4870
rect 3238 3576 3294 3632
rect 3974 3340 3976 3360
rect 3976 3340 4028 3360
rect 4028 3340 4030 3360
rect 3974 3304 4030 3340
rect 2870 1672 2926 1728
rect 4344 3834 4400 3836
rect 4424 3834 4480 3836
rect 4504 3834 4560 3836
rect 4584 3834 4640 3836
rect 4344 3782 4390 3834
rect 4390 3782 4400 3834
rect 4424 3782 4454 3834
rect 4454 3782 4466 3834
rect 4466 3782 4480 3834
rect 4504 3782 4518 3834
rect 4518 3782 4530 3834
rect 4530 3782 4560 3834
rect 4584 3782 4594 3834
rect 4594 3782 4640 3834
rect 4344 3780 4400 3782
rect 4424 3780 4480 3782
rect 4504 3780 4560 3782
rect 4584 3780 4640 3782
rect 4526 3576 4582 3632
rect 4344 2746 4400 2748
rect 4424 2746 4480 2748
rect 4504 2746 4560 2748
rect 4584 2746 4640 2748
rect 4344 2694 4390 2746
rect 4390 2694 4400 2746
rect 4424 2694 4454 2746
rect 4454 2694 4466 2746
rect 4466 2694 4480 2746
rect 4504 2694 4518 2746
rect 4518 2694 4530 2746
rect 4530 2694 4560 2746
rect 4584 2694 4594 2746
rect 4594 2694 4640 2746
rect 4344 2692 4400 2694
rect 4424 2692 4480 2694
rect 4504 2692 4560 2694
rect 4584 2692 4640 2694
rect 6182 14728 6238 14784
rect 6642 20460 6698 20496
rect 6642 20440 6644 20460
rect 6644 20440 6696 20460
rect 6696 20440 6698 20460
rect 6734 18708 6736 18728
rect 6736 18708 6788 18728
rect 6788 18708 6790 18728
rect 6734 18672 6790 18708
rect 6550 15952 6606 16008
rect 5998 12180 6000 12200
rect 6000 12180 6052 12200
rect 6052 12180 6054 12200
rect 5354 6568 5410 6624
rect 5998 12144 6054 12180
rect 6550 12144 6606 12200
rect 6642 10512 6698 10568
rect 7733 21786 7789 21788
rect 7813 21786 7869 21788
rect 7893 21786 7949 21788
rect 7973 21786 8029 21788
rect 7733 21734 7779 21786
rect 7779 21734 7789 21786
rect 7813 21734 7843 21786
rect 7843 21734 7855 21786
rect 7855 21734 7869 21786
rect 7893 21734 7907 21786
rect 7907 21734 7919 21786
rect 7919 21734 7949 21786
rect 7973 21734 7983 21786
rect 7983 21734 8029 21786
rect 7733 21732 7789 21734
rect 7813 21732 7869 21734
rect 7893 21732 7949 21734
rect 7973 21732 8029 21734
rect 7378 20576 7434 20632
rect 7733 20698 7789 20700
rect 7813 20698 7869 20700
rect 7893 20698 7949 20700
rect 7973 20698 8029 20700
rect 7733 20646 7779 20698
rect 7779 20646 7789 20698
rect 7813 20646 7843 20698
rect 7843 20646 7855 20698
rect 7855 20646 7869 20698
rect 7893 20646 7907 20698
rect 7907 20646 7919 20698
rect 7919 20646 7949 20698
rect 7973 20646 7983 20698
rect 7983 20646 8029 20698
rect 7733 20644 7789 20646
rect 7813 20644 7869 20646
rect 7893 20644 7949 20646
rect 7973 20644 8029 20646
rect 7562 19760 7618 19816
rect 7733 19610 7789 19612
rect 7813 19610 7869 19612
rect 7893 19610 7949 19612
rect 7973 19610 8029 19612
rect 7733 19558 7779 19610
rect 7779 19558 7789 19610
rect 7813 19558 7843 19610
rect 7843 19558 7855 19610
rect 7855 19558 7869 19610
rect 7893 19558 7907 19610
rect 7907 19558 7919 19610
rect 7919 19558 7949 19610
rect 7973 19558 7983 19610
rect 7983 19558 8029 19610
rect 7733 19556 7789 19558
rect 7813 19556 7869 19558
rect 7893 19556 7949 19558
rect 7973 19556 8029 19558
rect 7194 18708 7196 18728
rect 7196 18708 7248 18728
rect 7248 18708 7250 18728
rect 7194 18672 7250 18708
rect 7286 16532 7288 16552
rect 7288 16532 7340 16552
rect 7340 16532 7342 16552
rect 7286 16496 7342 16532
rect 7733 18522 7789 18524
rect 7813 18522 7869 18524
rect 7893 18522 7949 18524
rect 7973 18522 8029 18524
rect 7733 18470 7779 18522
rect 7779 18470 7789 18522
rect 7813 18470 7843 18522
rect 7843 18470 7855 18522
rect 7855 18470 7869 18522
rect 7893 18470 7907 18522
rect 7907 18470 7919 18522
rect 7919 18470 7949 18522
rect 7973 18470 7983 18522
rect 7983 18470 8029 18522
rect 7733 18468 7789 18470
rect 7813 18468 7869 18470
rect 7893 18468 7949 18470
rect 7973 18468 8029 18470
rect 7733 17434 7789 17436
rect 7813 17434 7869 17436
rect 7893 17434 7949 17436
rect 7973 17434 8029 17436
rect 7733 17382 7779 17434
rect 7779 17382 7789 17434
rect 7813 17382 7843 17434
rect 7843 17382 7855 17434
rect 7855 17382 7869 17434
rect 7893 17382 7907 17434
rect 7907 17382 7919 17434
rect 7919 17382 7949 17434
rect 7973 17382 7983 17434
rect 7983 17382 8029 17434
rect 7733 17380 7789 17382
rect 7813 17380 7869 17382
rect 7893 17380 7949 17382
rect 7973 17380 8029 17382
rect 8758 20460 8814 20496
rect 8758 20440 8760 20460
rect 8760 20440 8812 20460
rect 8812 20440 8814 20460
rect 8482 17620 8484 17640
rect 8484 17620 8536 17640
rect 8536 17620 8538 17640
rect 8482 17584 8538 17620
rect 7733 16346 7789 16348
rect 7813 16346 7869 16348
rect 7893 16346 7949 16348
rect 7973 16346 8029 16348
rect 7733 16294 7779 16346
rect 7779 16294 7789 16346
rect 7813 16294 7843 16346
rect 7843 16294 7855 16346
rect 7855 16294 7869 16346
rect 7893 16294 7907 16346
rect 7907 16294 7919 16346
rect 7919 16294 7949 16346
rect 7973 16294 7983 16346
rect 7983 16294 8029 16346
rect 7733 16292 7789 16294
rect 7813 16292 7869 16294
rect 7893 16292 7949 16294
rect 7973 16292 8029 16294
rect 7733 15258 7789 15260
rect 7813 15258 7869 15260
rect 7893 15258 7949 15260
rect 7973 15258 8029 15260
rect 7733 15206 7779 15258
rect 7779 15206 7789 15258
rect 7813 15206 7843 15258
rect 7843 15206 7855 15258
rect 7855 15206 7869 15258
rect 7893 15206 7907 15258
rect 7907 15206 7919 15258
rect 7919 15206 7949 15258
rect 7973 15206 7983 15258
rect 7983 15206 8029 15258
rect 7733 15204 7789 15206
rect 7813 15204 7869 15206
rect 7893 15204 7949 15206
rect 7973 15204 8029 15206
rect 6366 5752 6422 5808
rect 7194 9016 7250 9072
rect 7470 14048 7526 14104
rect 7746 15020 7802 15056
rect 7746 15000 7748 15020
rect 7748 15000 7800 15020
rect 7800 15000 7802 15020
rect 7733 14170 7789 14172
rect 7813 14170 7869 14172
rect 7893 14170 7949 14172
rect 7973 14170 8029 14172
rect 7733 14118 7779 14170
rect 7779 14118 7789 14170
rect 7813 14118 7843 14170
rect 7843 14118 7855 14170
rect 7855 14118 7869 14170
rect 7893 14118 7907 14170
rect 7907 14118 7919 14170
rect 7919 14118 7949 14170
rect 7973 14118 7983 14170
rect 7983 14118 8029 14170
rect 7733 14116 7789 14118
rect 7813 14116 7869 14118
rect 7893 14116 7949 14118
rect 7973 14116 8029 14118
rect 7733 13082 7789 13084
rect 7813 13082 7869 13084
rect 7893 13082 7949 13084
rect 7973 13082 8029 13084
rect 7733 13030 7779 13082
rect 7779 13030 7789 13082
rect 7813 13030 7843 13082
rect 7843 13030 7855 13082
rect 7855 13030 7869 13082
rect 7893 13030 7907 13082
rect 7907 13030 7919 13082
rect 7919 13030 7949 13082
rect 7973 13030 7983 13082
rect 7983 13030 8029 13082
rect 7733 13028 7789 13030
rect 7813 13028 7869 13030
rect 7893 13028 7949 13030
rect 7973 13028 8029 13030
rect 7378 9968 7434 10024
rect 7733 11994 7789 11996
rect 7813 11994 7869 11996
rect 7893 11994 7949 11996
rect 7973 11994 8029 11996
rect 7733 11942 7779 11994
rect 7779 11942 7789 11994
rect 7813 11942 7843 11994
rect 7843 11942 7855 11994
rect 7855 11942 7869 11994
rect 7893 11942 7907 11994
rect 7907 11942 7919 11994
rect 7919 11942 7949 11994
rect 7973 11942 7983 11994
rect 7983 11942 8029 11994
rect 7733 11940 7789 11942
rect 7813 11940 7869 11942
rect 7893 11940 7949 11942
rect 7973 11940 8029 11942
rect 7733 10906 7789 10908
rect 7813 10906 7869 10908
rect 7893 10906 7949 10908
rect 7973 10906 8029 10908
rect 7733 10854 7779 10906
rect 7779 10854 7789 10906
rect 7813 10854 7843 10906
rect 7843 10854 7855 10906
rect 7855 10854 7869 10906
rect 7893 10854 7907 10906
rect 7907 10854 7919 10906
rect 7919 10854 7949 10906
rect 7973 10854 7983 10906
rect 7983 10854 8029 10906
rect 7733 10852 7789 10854
rect 7813 10852 7869 10854
rect 7893 10852 7949 10854
rect 7973 10852 8029 10854
rect 7562 10512 7618 10568
rect 7286 6976 7342 7032
rect 7010 6160 7066 6216
rect 7102 4528 7158 4584
rect 7470 6296 7526 6352
rect 7470 6160 7526 6216
rect 8298 12144 8354 12200
rect 7733 9818 7789 9820
rect 7813 9818 7869 9820
rect 7893 9818 7949 9820
rect 7973 9818 8029 9820
rect 7733 9766 7779 9818
rect 7779 9766 7789 9818
rect 7813 9766 7843 9818
rect 7843 9766 7855 9818
rect 7855 9766 7869 9818
rect 7893 9766 7907 9818
rect 7907 9766 7919 9818
rect 7919 9766 7949 9818
rect 7973 9766 7983 9818
rect 7983 9766 8029 9818
rect 7733 9764 7789 9766
rect 7813 9764 7869 9766
rect 7893 9764 7949 9766
rect 7973 9764 8029 9766
rect 8114 9560 8170 9616
rect 7733 8730 7789 8732
rect 7813 8730 7869 8732
rect 7893 8730 7949 8732
rect 7973 8730 8029 8732
rect 7733 8678 7779 8730
rect 7779 8678 7789 8730
rect 7813 8678 7843 8730
rect 7843 8678 7855 8730
rect 7855 8678 7869 8730
rect 7893 8678 7907 8730
rect 7907 8678 7919 8730
rect 7919 8678 7949 8730
rect 7973 8678 7983 8730
rect 7983 8678 8029 8730
rect 7733 8676 7789 8678
rect 7813 8676 7869 8678
rect 7893 8676 7949 8678
rect 7973 8676 8029 8678
rect 7838 7948 7894 7984
rect 7838 7928 7840 7948
rect 7840 7928 7892 7948
rect 7892 7928 7894 7948
rect 7733 7642 7789 7644
rect 7813 7642 7869 7644
rect 7893 7642 7949 7644
rect 7973 7642 8029 7644
rect 7733 7590 7779 7642
rect 7779 7590 7789 7642
rect 7813 7590 7843 7642
rect 7843 7590 7855 7642
rect 7855 7590 7869 7642
rect 7893 7590 7907 7642
rect 7907 7590 7919 7642
rect 7919 7590 7949 7642
rect 7973 7590 7983 7642
rect 7983 7590 8029 7642
rect 7733 7588 7789 7590
rect 7813 7588 7869 7590
rect 7893 7588 7949 7590
rect 7973 7588 8029 7590
rect 8298 10260 8354 10296
rect 8298 10240 8300 10260
rect 8300 10240 8352 10260
rect 8352 10240 8354 10260
rect 8298 7404 8354 7440
rect 8298 7384 8300 7404
rect 8300 7384 8352 7404
rect 8352 7384 8354 7404
rect 7733 6554 7789 6556
rect 7813 6554 7869 6556
rect 7893 6554 7949 6556
rect 7973 6554 8029 6556
rect 7733 6502 7779 6554
rect 7779 6502 7789 6554
rect 7813 6502 7843 6554
rect 7843 6502 7855 6554
rect 7855 6502 7869 6554
rect 7893 6502 7907 6554
rect 7907 6502 7919 6554
rect 7919 6502 7949 6554
rect 7973 6502 7983 6554
rect 7983 6502 8029 6554
rect 7733 6500 7789 6502
rect 7813 6500 7869 6502
rect 7893 6500 7949 6502
rect 7973 6500 8029 6502
rect 7733 5466 7789 5468
rect 7813 5466 7869 5468
rect 7893 5466 7949 5468
rect 7973 5466 8029 5468
rect 7733 5414 7779 5466
rect 7779 5414 7789 5466
rect 7813 5414 7843 5466
rect 7843 5414 7855 5466
rect 7855 5414 7869 5466
rect 7893 5414 7907 5466
rect 7907 5414 7919 5466
rect 7919 5414 7949 5466
rect 7973 5414 7983 5466
rect 7983 5414 8029 5466
rect 7733 5412 7789 5414
rect 7813 5412 7869 5414
rect 7893 5412 7949 5414
rect 7973 5412 8029 5414
rect 7733 4378 7789 4380
rect 7813 4378 7869 4380
rect 7893 4378 7949 4380
rect 7973 4378 8029 4380
rect 7733 4326 7779 4378
rect 7779 4326 7789 4378
rect 7813 4326 7843 4378
rect 7843 4326 7855 4378
rect 7855 4326 7869 4378
rect 7893 4326 7907 4378
rect 7907 4326 7919 4378
rect 7919 4326 7949 4378
rect 7973 4326 7983 4378
rect 7983 4326 8029 4378
rect 7733 4324 7789 4326
rect 7813 4324 7869 4326
rect 7893 4324 7949 4326
rect 7973 4324 8029 4326
rect 7733 3290 7789 3292
rect 7813 3290 7869 3292
rect 7893 3290 7949 3292
rect 7973 3290 8029 3292
rect 7733 3238 7779 3290
rect 7779 3238 7789 3290
rect 7813 3238 7843 3290
rect 7843 3238 7855 3290
rect 7855 3238 7869 3290
rect 7893 3238 7907 3290
rect 7907 3238 7919 3290
rect 7919 3238 7949 3290
rect 7973 3238 7983 3290
rect 7983 3238 8029 3290
rect 7733 3236 7789 3238
rect 7813 3236 7869 3238
rect 7893 3236 7949 3238
rect 7973 3236 8029 3238
rect 7733 2202 7789 2204
rect 7813 2202 7869 2204
rect 7893 2202 7949 2204
rect 7973 2202 8029 2204
rect 7733 2150 7779 2202
rect 7779 2150 7789 2202
rect 7813 2150 7843 2202
rect 7843 2150 7855 2202
rect 7855 2150 7869 2202
rect 7893 2150 7907 2202
rect 7907 2150 7919 2202
rect 7919 2150 7949 2202
rect 7973 2150 7983 2202
rect 7983 2150 8029 2202
rect 7733 2148 7789 2150
rect 7813 2148 7869 2150
rect 7893 2148 7949 2150
rect 7973 2148 8029 2150
rect 8850 17176 8906 17232
rect 8850 12960 8906 13016
rect 11122 22330 11178 22332
rect 11202 22330 11258 22332
rect 11282 22330 11338 22332
rect 11362 22330 11418 22332
rect 11122 22278 11168 22330
rect 11168 22278 11178 22330
rect 11202 22278 11232 22330
rect 11232 22278 11244 22330
rect 11244 22278 11258 22330
rect 11282 22278 11296 22330
rect 11296 22278 11308 22330
rect 11308 22278 11338 22330
rect 11362 22278 11372 22330
rect 11372 22278 11418 22330
rect 11122 22276 11178 22278
rect 11202 22276 11258 22278
rect 11282 22276 11338 22278
rect 11362 22276 11418 22278
rect 10046 21392 10102 21448
rect 9310 19372 9366 19408
rect 9310 19352 9312 19372
rect 9312 19352 9364 19372
rect 9364 19352 9366 19372
rect 9310 16496 9366 16552
rect 9310 14864 9366 14920
rect 10138 20984 10194 21040
rect 10046 20748 10048 20768
rect 10048 20748 10100 20768
rect 10100 20748 10102 20768
rect 10046 20712 10102 20748
rect 9770 19488 9826 19544
rect 9494 14592 9550 14648
rect 9218 14048 9274 14104
rect 9494 14048 9550 14104
rect 9126 12588 9128 12608
rect 9128 12588 9180 12608
rect 9180 12588 9182 12608
rect 9126 12552 9182 12588
rect 9126 12416 9182 12472
rect 8942 9696 8998 9752
rect 9678 14456 9734 14512
rect 10230 17720 10286 17776
rect 10230 16652 10286 16688
rect 10230 16632 10232 16652
rect 10232 16632 10284 16652
rect 10284 16632 10286 16652
rect 10230 15952 10286 16008
rect 9954 13912 10010 13968
rect 10138 13404 10140 13424
rect 10140 13404 10192 13424
rect 10192 13404 10194 13424
rect 10138 13368 10194 13404
rect 9402 12552 9458 12608
rect 9494 12280 9550 12336
rect 9126 6840 9182 6896
rect 9862 12688 9918 12744
rect 9034 5480 9090 5536
rect 9310 5208 9366 5264
rect 9218 4800 9274 4856
rect 9494 9968 9550 10024
rect 9494 9716 9550 9752
rect 9494 9696 9496 9716
rect 9496 9696 9548 9716
rect 9548 9696 9550 9716
rect 9494 5480 9550 5536
rect 9586 5344 9642 5400
rect 9586 5092 9642 5128
rect 9586 5072 9588 5092
rect 9588 5072 9640 5092
rect 9640 5072 9642 5092
rect 9586 4820 9642 4856
rect 9586 4800 9588 4820
rect 9588 4800 9640 4820
rect 9640 4800 9642 4820
rect 9954 10240 10010 10296
rect 9954 7520 10010 7576
rect 9862 5108 9864 5128
rect 9864 5108 9916 5128
rect 9916 5108 9918 5128
rect 9862 5072 9918 5108
rect 10322 12144 10378 12200
rect 10414 10260 10470 10296
rect 10414 10240 10416 10260
rect 10416 10240 10468 10260
rect 10468 10240 10470 10260
rect 11122 21242 11178 21244
rect 11202 21242 11258 21244
rect 11282 21242 11338 21244
rect 11362 21242 11418 21244
rect 11122 21190 11168 21242
rect 11168 21190 11178 21242
rect 11202 21190 11232 21242
rect 11232 21190 11244 21242
rect 11244 21190 11258 21242
rect 11282 21190 11296 21242
rect 11296 21190 11308 21242
rect 11308 21190 11338 21242
rect 11362 21190 11372 21242
rect 11372 21190 11418 21242
rect 11122 21188 11178 21190
rect 11202 21188 11258 21190
rect 11282 21188 11338 21190
rect 11362 21188 11418 21190
rect 11058 21004 11114 21040
rect 11058 20984 11060 21004
rect 11060 20984 11112 21004
rect 11112 20984 11114 21004
rect 10782 20848 10838 20904
rect 11122 20154 11178 20156
rect 11202 20154 11258 20156
rect 11282 20154 11338 20156
rect 11362 20154 11418 20156
rect 11122 20102 11168 20154
rect 11168 20102 11178 20154
rect 11202 20102 11232 20154
rect 11232 20102 11244 20154
rect 11244 20102 11258 20154
rect 11282 20102 11296 20154
rect 11296 20102 11308 20154
rect 11308 20102 11338 20154
rect 11362 20102 11372 20154
rect 11372 20102 11418 20154
rect 11122 20100 11178 20102
rect 11202 20100 11258 20102
rect 11282 20100 11338 20102
rect 11362 20100 11418 20102
rect 11518 20032 11574 20088
rect 12070 20984 12126 21040
rect 12070 20748 12072 20768
rect 12072 20748 12124 20768
rect 12124 20748 12126 20768
rect 12070 20712 12126 20748
rect 11122 19066 11178 19068
rect 11202 19066 11258 19068
rect 11282 19066 11338 19068
rect 11362 19066 11418 19068
rect 11122 19014 11168 19066
rect 11168 19014 11178 19066
rect 11202 19014 11232 19066
rect 11232 19014 11244 19066
rect 11244 19014 11258 19066
rect 11282 19014 11296 19066
rect 11296 19014 11308 19066
rect 11308 19014 11338 19066
rect 11362 19014 11372 19066
rect 11372 19014 11418 19066
rect 11122 19012 11178 19014
rect 11202 19012 11258 19014
rect 11282 19012 11338 19014
rect 11362 19012 11418 19014
rect 10782 18828 10838 18864
rect 10782 18808 10784 18828
rect 10784 18808 10836 18828
rect 10836 18808 10838 18828
rect 10782 17176 10838 17232
rect 11122 17978 11178 17980
rect 11202 17978 11258 17980
rect 11282 17978 11338 17980
rect 11362 17978 11418 17980
rect 11122 17926 11168 17978
rect 11168 17926 11178 17978
rect 11202 17926 11232 17978
rect 11232 17926 11244 17978
rect 11244 17926 11258 17978
rect 11282 17926 11296 17978
rect 11296 17926 11308 17978
rect 11308 17926 11338 17978
rect 11362 17926 11372 17978
rect 11372 17926 11418 17978
rect 11122 17924 11178 17926
rect 11202 17924 11258 17926
rect 11282 17924 11338 17926
rect 11362 17924 11418 17926
rect 11518 17584 11574 17640
rect 11122 16890 11178 16892
rect 11202 16890 11258 16892
rect 11282 16890 11338 16892
rect 11362 16890 11418 16892
rect 11122 16838 11168 16890
rect 11168 16838 11178 16890
rect 11202 16838 11232 16890
rect 11232 16838 11244 16890
rect 11244 16838 11258 16890
rect 11282 16838 11296 16890
rect 11296 16838 11308 16890
rect 11308 16838 11338 16890
rect 11362 16838 11372 16890
rect 11372 16838 11418 16890
rect 11122 16836 11178 16838
rect 11202 16836 11258 16838
rect 11282 16836 11338 16838
rect 11362 16836 11418 16838
rect 10690 14864 10746 14920
rect 10598 14456 10654 14512
rect 11122 15802 11178 15804
rect 11202 15802 11258 15804
rect 11282 15802 11338 15804
rect 11362 15802 11418 15804
rect 11122 15750 11168 15802
rect 11168 15750 11178 15802
rect 11202 15750 11232 15802
rect 11232 15750 11244 15802
rect 11244 15750 11258 15802
rect 11282 15750 11296 15802
rect 11296 15750 11308 15802
rect 11308 15750 11338 15802
rect 11362 15750 11372 15802
rect 11372 15750 11418 15802
rect 11122 15748 11178 15750
rect 11202 15748 11258 15750
rect 11282 15748 11338 15750
rect 11362 15748 11418 15750
rect 11886 19352 11942 19408
rect 11886 18264 11942 18320
rect 11978 17312 12034 17368
rect 11978 16496 12034 16552
rect 10966 14728 11022 14784
rect 11122 14714 11178 14716
rect 11202 14714 11258 14716
rect 11282 14714 11338 14716
rect 11362 14714 11418 14716
rect 11122 14662 11168 14714
rect 11168 14662 11178 14714
rect 11202 14662 11232 14714
rect 11232 14662 11244 14714
rect 11244 14662 11258 14714
rect 11282 14662 11296 14714
rect 11296 14662 11308 14714
rect 11308 14662 11338 14714
rect 11362 14662 11372 14714
rect 11372 14662 11418 14714
rect 11122 14660 11178 14662
rect 11202 14660 11258 14662
rect 11282 14660 11338 14662
rect 11362 14660 11418 14662
rect 11122 13626 11178 13628
rect 11202 13626 11258 13628
rect 11282 13626 11338 13628
rect 11362 13626 11418 13628
rect 11122 13574 11168 13626
rect 11168 13574 11178 13626
rect 11202 13574 11232 13626
rect 11232 13574 11244 13626
rect 11244 13574 11258 13626
rect 11282 13574 11296 13626
rect 11296 13574 11308 13626
rect 11308 13574 11338 13626
rect 11362 13574 11372 13626
rect 11372 13574 11418 13626
rect 11122 13572 11178 13574
rect 11202 13572 11258 13574
rect 11282 13572 11338 13574
rect 11362 13572 11418 13574
rect 11122 12538 11178 12540
rect 11202 12538 11258 12540
rect 11282 12538 11338 12540
rect 11362 12538 11418 12540
rect 11122 12486 11168 12538
rect 11168 12486 11178 12538
rect 11202 12486 11232 12538
rect 11232 12486 11244 12538
rect 11244 12486 11258 12538
rect 11282 12486 11296 12538
rect 11296 12486 11308 12538
rect 11308 12486 11338 12538
rect 11362 12486 11372 12538
rect 11372 12486 11418 12538
rect 11122 12484 11178 12486
rect 11202 12484 11258 12486
rect 11282 12484 11338 12486
rect 11362 12484 11418 12486
rect 10506 9560 10562 9616
rect 9678 3596 9734 3632
rect 9678 3576 9680 3596
rect 9680 3576 9732 3596
rect 9732 3576 9734 3596
rect 11122 11450 11178 11452
rect 11202 11450 11258 11452
rect 11282 11450 11338 11452
rect 11362 11450 11418 11452
rect 11122 11398 11168 11450
rect 11168 11398 11178 11450
rect 11202 11398 11232 11450
rect 11232 11398 11244 11450
rect 11244 11398 11258 11450
rect 11282 11398 11296 11450
rect 11296 11398 11308 11450
rect 11308 11398 11338 11450
rect 11362 11398 11372 11450
rect 11372 11398 11418 11450
rect 11122 11396 11178 11398
rect 11202 11396 11258 11398
rect 11282 11396 11338 11398
rect 11362 11396 11418 11398
rect 11702 12280 11758 12336
rect 11122 10362 11178 10364
rect 11202 10362 11258 10364
rect 11282 10362 11338 10364
rect 11362 10362 11418 10364
rect 11122 10310 11168 10362
rect 11168 10310 11178 10362
rect 11202 10310 11232 10362
rect 11232 10310 11244 10362
rect 11244 10310 11258 10362
rect 11282 10310 11296 10362
rect 11296 10310 11308 10362
rect 11308 10310 11338 10362
rect 11362 10310 11372 10362
rect 11372 10310 11418 10362
rect 11122 10308 11178 10310
rect 11202 10308 11258 10310
rect 11282 10308 11338 10310
rect 11362 10308 11418 10310
rect 11122 9274 11178 9276
rect 11202 9274 11258 9276
rect 11282 9274 11338 9276
rect 11362 9274 11418 9276
rect 11122 9222 11168 9274
rect 11168 9222 11178 9274
rect 11202 9222 11232 9274
rect 11232 9222 11244 9274
rect 11244 9222 11258 9274
rect 11282 9222 11296 9274
rect 11296 9222 11308 9274
rect 11308 9222 11338 9274
rect 11362 9222 11372 9274
rect 11372 9222 11418 9274
rect 11122 9220 11178 9222
rect 11202 9220 11258 9222
rect 11282 9220 11338 9222
rect 11362 9220 11418 9222
rect 10966 8880 11022 8936
rect 11122 8186 11178 8188
rect 11202 8186 11258 8188
rect 11282 8186 11338 8188
rect 11362 8186 11418 8188
rect 11122 8134 11168 8186
rect 11168 8134 11178 8186
rect 11202 8134 11232 8186
rect 11232 8134 11244 8186
rect 11244 8134 11258 8186
rect 11282 8134 11296 8186
rect 11296 8134 11308 8186
rect 11308 8134 11338 8186
rect 11362 8134 11372 8186
rect 11372 8134 11418 8186
rect 11122 8132 11178 8134
rect 11202 8132 11258 8134
rect 11282 8132 11338 8134
rect 11362 8132 11418 8134
rect 11242 7928 11298 7984
rect 11150 7248 11206 7304
rect 11122 7098 11178 7100
rect 11202 7098 11258 7100
rect 11282 7098 11338 7100
rect 11362 7098 11418 7100
rect 11122 7046 11168 7098
rect 11168 7046 11178 7098
rect 11202 7046 11232 7098
rect 11232 7046 11244 7098
rect 11244 7046 11258 7098
rect 11282 7046 11296 7098
rect 11296 7046 11308 7098
rect 11308 7046 11338 7098
rect 11362 7046 11372 7098
rect 11372 7046 11418 7098
rect 11122 7044 11178 7046
rect 11202 7044 11258 7046
rect 11282 7044 11338 7046
rect 11362 7044 11418 7046
rect 11122 6010 11178 6012
rect 11202 6010 11258 6012
rect 11282 6010 11338 6012
rect 11362 6010 11418 6012
rect 11122 5958 11168 6010
rect 11168 5958 11178 6010
rect 11202 5958 11232 6010
rect 11232 5958 11244 6010
rect 11244 5958 11258 6010
rect 11282 5958 11296 6010
rect 11296 5958 11308 6010
rect 11308 5958 11338 6010
rect 11362 5958 11372 6010
rect 11372 5958 11418 6010
rect 11122 5956 11178 5958
rect 11202 5956 11258 5958
rect 11282 5956 11338 5958
rect 11362 5956 11418 5958
rect 11702 7812 11758 7848
rect 11702 7792 11704 7812
rect 11704 7792 11756 7812
rect 11756 7792 11758 7812
rect 11610 6568 11666 6624
rect 11122 4922 11178 4924
rect 11202 4922 11258 4924
rect 11282 4922 11338 4924
rect 11362 4922 11418 4924
rect 11122 4870 11168 4922
rect 11168 4870 11178 4922
rect 11202 4870 11232 4922
rect 11232 4870 11244 4922
rect 11244 4870 11258 4922
rect 11282 4870 11296 4922
rect 11296 4870 11308 4922
rect 11308 4870 11338 4922
rect 11362 4870 11372 4922
rect 11372 4870 11418 4922
rect 11122 4868 11178 4870
rect 11202 4868 11258 4870
rect 11282 4868 11338 4870
rect 11362 4868 11418 4870
rect 11122 3834 11178 3836
rect 11202 3834 11258 3836
rect 11282 3834 11338 3836
rect 11362 3834 11418 3836
rect 11122 3782 11168 3834
rect 11168 3782 11178 3834
rect 11202 3782 11232 3834
rect 11232 3782 11244 3834
rect 11244 3782 11258 3834
rect 11282 3782 11296 3834
rect 11296 3782 11308 3834
rect 11308 3782 11338 3834
rect 11362 3782 11372 3834
rect 11372 3782 11418 3834
rect 11122 3780 11178 3782
rect 11202 3780 11258 3782
rect 11282 3780 11338 3782
rect 11362 3780 11418 3782
rect 11122 2746 11178 2748
rect 11202 2746 11258 2748
rect 11282 2746 11338 2748
rect 11362 2746 11418 2748
rect 11122 2694 11168 2746
rect 11168 2694 11178 2746
rect 11202 2694 11232 2746
rect 11232 2694 11244 2746
rect 11244 2694 11258 2746
rect 11282 2694 11296 2746
rect 11296 2694 11308 2746
rect 11308 2694 11338 2746
rect 11362 2694 11372 2746
rect 11372 2694 11418 2746
rect 11122 2692 11178 2694
rect 11202 2692 11258 2694
rect 11282 2692 11338 2694
rect 11362 2692 11418 2694
rect 11978 9460 11980 9480
rect 11980 9460 12032 9480
rect 12032 9460 12034 9480
rect 11978 9424 12034 9460
rect 12346 19488 12402 19544
rect 12530 18808 12586 18864
rect 12898 20032 12954 20088
rect 12806 19388 12808 19408
rect 12808 19388 12860 19408
rect 12860 19388 12862 19408
rect 12806 19352 12862 19388
rect 12346 17856 12402 17912
rect 12346 17040 12402 17096
rect 13174 18828 13230 18864
rect 13174 18808 13176 18828
rect 13176 18808 13228 18828
rect 13228 18808 13230 18828
rect 12806 17040 12862 17096
rect 12346 12960 12402 13016
rect 12622 13368 12678 13424
rect 12438 12436 12494 12472
rect 12438 12416 12440 12436
rect 12440 12416 12492 12436
rect 12492 12416 12494 12436
rect 12254 11736 12310 11792
rect 12530 11736 12586 11792
rect 12990 11500 12992 11520
rect 12992 11500 13044 11520
rect 13044 11500 13046 11520
rect 12990 11464 13046 11500
rect 12254 7540 12310 7576
rect 12254 7520 12256 7540
rect 12256 7520 12308 7540
rect 12308 7520 12310 7540
rect 13082 10376 13138 10432
rect 12806 9424 12862 9480
rect 12622 7520 12678 7576
rect 12806 8472 12862 8528
rect 12346 6568 12402 6624
rect 12898 5072 12954 5128
rect 12438 3188 12494 3224
rect 12438 3168 12440 3188
rect 12440 3168 12492 3188
rect 12492 3168 12494 3188
rect 12898 3168 12954 3224
rect 13726 19508 13782 19544
rect 13726 19488 13728 19508
rect 13728 19488 13780 19508
rect 13780 19488 13782 19508
rect 13542 17312 13598 17368
rect 13726 17040 13782 17096
rect 14510 21786 14566 21788
rect 14590 21786 14646 21788
rect 14670 21786 14726 21788
rect 14750 21786 14806 21788
rect 14510 21734 14556 21786
rect 14556 21734 14566 21786
rect 14590 21734 14620 21786
rect 14620 21734 14632 21786
rect 14632 21734 14646 21786
rect 14670 21734 14684 21786
rect 14684 21734 14696 21786
rect 14696 21734 14726 21786
rect 14750 21734 14760 21786
rect 14760 21734 14806 21786
rect 14510 21732 14566 21734
rect 14590 21732 14646 21734
rect 14670 21732 14726 21734
rect 14750 21732 14806 21734
rect 14370 21392 14426 21448
rect 14510 20698 14566 20700
rect 14590 20698 14646 20700
rect 14670 20698 14726 20700
rect 14750 20698 14806 20700
rect 14510 20646 14556 20698
rect 14556 20646 14566 20698
rect 14590 20646 14620 20698
rect 14620 20646 14632 20698
rect 14632 20646 14646 20698
rect 14670 20646 14684 20698
rect 14684 20646 14696 20698
rect 14696 20646 14726 20698
rect 14750 20646 14760 20698
rect 14760 20646 14806 20698
rect 14510 20644 14566 20646
rect 14590 20644 14646 20646
rect 14670 20644 14726 20646
rect 14750 20644 14806 20646
rect 14510 19610 14566 19612
rect 14590 19610 14646 19612
rect 14670 19610 14726 19612
rect 14750 19610 14806 19612
rect 14510 19558 14556 19610
rect 14556 19558 14566 19610
rect 14590 19558 14620 19610
rect 14620 19558 14632 19610
rect 14632 19558 14646 19610
rect 14670 19558 14684 19610
rect 14684 19558 14696 19610
rect 14696 19558 14726 19610
rect 14750 19558 14760 19610
rect 14760 19558 14806 19610
rect 14510 19556 14566 19558
rect 14590 19556 14646 19558
rect 14670 19556 14726 19558
rect 14750 19556 14806 19558
rect 14510 18522 14566 18524
rect 14590 18522 14646 18524
rect 14670 18522 14726 18524
rect 14750 18522 14806 18524
rect 14510 18470 14556 18522
rect 14556 18470 14566 18522
rect 14590 18470 14620 18522
rect 14620 18470 14632 18522
rect 14632 18470 14646 18522
rect 14670 18470 14684 18522
rect 14684 18470 14696 18522
rect 14696 18470 14726 18522
rect 14750 18470 14760 18522
rect 14760 18470 14806 18522
rect 14510 18468 14566 18470
rect 14590 18468 14646 18470
rect 14670 18468 14726 18470
rect 14750 18468 14806 18470
rect 14922 19216 14978 19272
rect 14510 17434 14566 17436
rect 14590 17434 14646 17436
rect 14670 17434 14726 17436
rect 14750 17434 14806 17436
rect 14510 17382 14556 17434
rect 14556 17382 14566 17434
rect 14590 17382 14620 17434
rect 14620 17382 14632 17434
rect 14632 17382 14646 17434
rect 14670 17382 14684 17434
rect 14684 17382 14696 17434
rect 14696 17382 14726 17434
rect 14750 17382 14760 17434
rect 14760 17382 14806 17434
rect 14510 17380 14566 17382
rect 14590 17380 14646 17382
rect 14670 17380 14726 17382
rect 14750 17380 14806 17382
rect 14186 16788 14242 16824
rect 14186 16768 14188 16788
rect 14188 16768 14240 16788
rect 14240 16768 14242 16788
rect 14830 16768 14886 16824
rect 15474 17856 15530 17912
rect 14510 16346 14566 16348
rect 14590 16346 14646 16348
rect 14670 16346 14726 16348
rect 14750 16346 14806 16348
rect 14510 16294 14556 16346
rect 14556 16294 14566 16346
rect 14590 16294 14620 16346
rect 14620 16294 14632 16346
rect 14632 16294 14646 16346
rect 14670 16294 14684 16346
rect 14684 16294 14696 16346
rect 14696 16294 14726 16346
rect 14750 16294 14760 16346
rect 14760 16294 14806 16346
rect 14510 16292 14566 16294
rect 14590 16292 14646 16294
rect 14670 16292 14726 16294
rect 14750 16292 14806 16294
rect 14510 15258 14566 15260
rect 14590 15258 14646 15260
rect 14670 15258 14726 15260
rect 14750 15258 14806 15260
rect 14510 15206 14556 15258
rect 14556 15206 14566 15258
rect 14590 15206 14620 15258
rect 14620 15206 14632 15258
rect 14632 15206 14646 15258
rect 14670 15206 14684 15258
rect 14684 15206 14696 15258
rect 14696 15206 14726 15258
rect 14750 15206 14760 15258
rect 14760 15206 14806 15258
rect 14510 15204 14566 15206
rect 14590 15204 14646 15206
rect 14670 15204 14726 15206
rect 14750 15204 14806 15206
rect 14738 14476 14794 14512
rect 14738 14456 14740 14476
rect 14740 14456 14792 14476
rect 14792 14456 14794 14476
rect 14510 14170 14566 14172
rect 14590 14170 14646 14172
rect 14670 14170 14726 14172
rect 14750 14170 14806 14172
rect 14510 14118 14556 14170
rect 14556 14118 14566 14170
rect 14590 14118 14620 14170
rect 14620 14118 14632 14170
rect 14632 14118 14646 14170
rect 14670 14118 14684 14170
rect 14684 14118 14696 14170
rect 14696 14118 14726 14170
rect 14750 14118 14760 14170
rect 14760 14118 14806 14170
rect 14510 14116 14566 14118
rect 14590 14116 14646 14118
rect 14670 14116 14726 14118
rect 14750 14116 14806 14118
rect 14510 13082 14566 13084
rect 14590 13082 14646 13084
rect 14670 13082 14726 13084
rect 14750 13082 14806 13084
rect 14510 13030 14556 13082
rect 14556 13030 14566 13082
rect 14590 13030 14620 13082
rect 14620 13030 14632 13082
rect 14632 13030 14646 13082
rect 14670 13030 14684 13082
rect 14684 13030 14696 13082
rect 14696 13030 14726 13082
rect 14750 13030 14760 13082
rect 14760 13030 14806 13082
rect 14510 13028 14566 13030
rect 14590 13028 14646 13030
rect 14670 13028 14726 13030
rect 14750 13028 14806 13030
rect 14462 12588 14464 12608
rect 14464 12588 14516 12608
rect 14516 12588 14518 12608
rect 14462 12552 14518 12588
rect 14554 12416 14610 12472
rect 14510 11994 14566 11996
rect 14590 11994 14646 11996
rect 14670 11994 14726 11996
rect 14750 11994 14806 11996
rect 14510 11942 14556 11994
rect 14556 11942 14566 11994
rect 14590 11942 14620 11994
rect 14620 11942 14632 11994
rect 14632 11942 14646 11994
rect 14670 11942 14684 11994
rect 14684 11942 14696 11994
rect 14696 11942 14726 11994
rect 14750 11942 14760 11994
rect 14760 11942 14806 11994
rect 14510 11940 14566 11942
rect 14590 11940 14646 11942
rect 14670 11940 14726 11942
rect 14750 11940 14806 11942
rect 14830 11348 14886 11384
rect 14830 11328 14832 11348
rect 14832 11328 14884 11348
rect 14884 11328 14886 11348
rect 14510 10906 14566 10908
rect 14590 10906 14646 10908
rect 14670 10906 14726 10908
rect 14750 10906 14806 10908
rect 14510 10854 14556 10906
rect 14556 10854 14566 10906
rect 14590 10854 14620 10906
rect 14620 10854 14632 10906
rect 14632 10854 14646 10906
rect 14670 10854 14684 10906
rect 14684 10854 14696 10906
rect 14696 10854 14726 10906
rect 14750 10854 14760 10906
rect 14760 10854 14806 10906
rect 14510 10852 14566 10854
rect 14590 10852 14646 10854
rect 14670 10852 14726 10854
rect 14750 10852 14806 10854
rect 13910 7520 13966 7576
rect 14510 9818 14566 9820
rect 14590 9818 14646 9820
rect 14670 9818 14726 9820
rect 14750 9818 14806 9820
rect 14510 9766 14556 9818
rect 14556 9766 14566 9818
rect 14590 9766 14620 9818
rect 14620 9766 14632 9818
rect 14632 9766 14646 9818
rect 14670 9766 14684 9818
rect 14684 9766 14696 9818
rect 14696 9766 14726 9818
rect 14750 9766 14760 9818
rect 14760 9766 14806 9818
rect 14510 9764 14566 9766
rect 14590 9764 14646 9766
rect 14670 9764 14726 9766
rect 14750 9764 14806 9766
rect 14510 8730 14566 8732
rect 14590 8730 14646 8732
rect 14670 8730 14726 8732
rect 14750 8730 14806 8732
rect 14510 8678 14556 8730
rect 14556 8678 14566 8730
rect 14590 8678 14620 8730
rect 14620 8678 14632 8730
rect 14632 8678 14646 8730
rect 14670 8678 14684 8730
rect 14684 8678 14696 8730
rect 14696 8678 14726 8730
rect 14750 8678 14760 8730
rect 14760 8678 14806 8730
rect 14510 8676 14566 8678
rect 14590 8676 14646 8678
rect 14670 8676 14726 8678
rect 14750 8676 14806 8678
rect 15106 13368 15162 13424
rect 15198 12552 15254 12608
rect 16486 20984 16542 21040
rect 16762 20984 16818 21040
rect 15750 15952 15806 16008
rect 15474 13268 15476 13288
rect 15476 13268 15528 13288
rect 15528 13268 15530 13288
rect 15474 13232 15530 13268
rect 15750 13776 15806 13832
rect 15658 13232 15714 13288
rect 15290 11328 15346 11384
rect 14370 8200 14426 8256
rect 14510 7642 14566 7644
rect 14590 7642 14646 7644
rect 14670 7642 14726 7644
rect 14750 7642 14806 7644
rect 14510 7590 14556 7642
rect 14556 7590 14566 7642
rect 14590 7590 14620 7642
rect 14620 7590 14632 7642
rect 14632 7590 14646 7642
rect 14670 7590 14684 7642
rect 14684 7590 14696 7642
rect 14696 7590 14726 7642
rect 14750 7590 14760 7642
rect 14760 7590 14806 7642
rect 14510 7588 14566 7590
rect 14590 7588 14646 7590
rect 14670 7588 14726 7590
rect 14750 7588 14806 7590
rect 14922 7928 14978 7984
rect 15106 8356 15162 8392
rect 15106 8336 15108 8356
rect 15108 8336 15160 8356
rect 15160 8336 15162 8356
rect 13818 5108 13820 5128
rect 13820 5108 13872 5128
rect 13872 5108 13874 5128
rect 13818 5072 13874 5108
rect 14510 6554 14566 6556
rect 14590 6554 14646 6556
rect 14670 6554 14726 6556
rect 14750 6554 14806 6556
rect 14510 6502 14556 6554
rect 14556 6502 14566 6554
rect 14590 6502 14620 6554
rect 14620 6502 14632 6554
rect 14632 6502 14646 6554
rect 14670 6502 14684 6554
rect 14684 6502 14696 6554
rect 14696 6502 14726 6554
rect 14750 6502 14760 6554
rect 14760 6502 14806 6554
rect 14510 6500 14566 6502
rect 14590 6500 14646 6502
rect 14670 6500 14726 6502
rect 14750 6500 14806 6502
rect 14510 5466 14566 5468
rect 14590 5466 14646 5468
rect 14670 5466 14726 5468
rect 14750 5466 14806 5468
rect 14510 5414 14556 5466
rect 14556 5414 14566 5466
rect 14590 5414 14620 5466
rect 14620 5414 14632 5466
rect 14632 5414 14646 5466
rect 14670 5414 14684 5466
rect 14684 5414 14696 5466
rect 14696 5414 14726 5466
rect 14750 5414 14760 5466
rect 14760 5414 14806 5466
rect 14510 5412 14566 5414
rect 14590 5412 14646 5414
rect 14670 5412 14726 5414
rect 14750 5412 14806 5414
rect 14738 5228 14794 5264
rect 14738 5208 14740 5228
rect 14740 5208 14792 5228
rect 14792 5208 14794 5228
rect 13910 3612 13912 3632
rect 13912 3612 13964 3632
rect 13964 3612 13966 3632
rect 13910 3576 13966 3612
rect 14510 4378 14566 4380
rect 14590 4378 14646 4380
rect 14670 4378 14726 4380
rect 14750 4378 14806 4380
rect 14510 4326 14556 4378
rect 14556 4326 14566 4378
rect 14590 4326 14620 4378
rect 14620 4326 14632 4378
rect 14632 4326 14646 4378
rect 14670 4326 14684 4378
rect 14684 4326 14696 4378
rect 14696 4326 14726 4378
rect 14750 4326 14760 4378
rect 14760 4326 14806 4378
rect 14510 4324 14566 4326
rect 14590 4324 14646 4326
rect 14670 4324 14726 4326
rect 14750 4324 14806 4326
rect 15382 6704 15438 6760
rect 14510 3290 14566 3292
rect 14590 3290 14646 3292
rect 14670 3290 14726 3292
rect 14750 3290 14806 3292
rect 14510 3238 14556 3290
rect 14556 3238 14566 3290
rect 14590 3238 14620 3290
rect 14620 3238 14632 3290
rect 14632 3238 14646 3290
rect 14670 3238 14684 3290
rect 14684 3238 14696 3290
rect 14696 3238 14726 3290
rect 14750 3238 14760 3290
rect 14760 3238 14806 3290
rect 14510 3236 14566 3238
rect 14590 3236 14646 3238
rect 14670 3236 14726 3238
rect 14750 3236 14806 3238
rect 15382 3304 15438 3360
rect 16118 14864 16174 14920
rect 15658 8880 15714 8936
rect 16026 11464 16082 11520
rect 16578 18284 16634 18320
rect 16578 18264 16580 18284
rect 16580 18264 16632 18284
rect 16632 18264 16634 18284
rect 16578 16632 16634 16688
rect 16394 15000 16450 15056
rect 17899 22330 17955 22332
rect 17979 22330 18035 22332
rect 18059 22330 18115 22332
rect 18139 22330 18195 22332
rect 17899 22278 17945 22330
rect 17945 22278 17955 22330
rect 17979 22278 18009 22330
rect 18009 22278 18021 22330
rect 18021 22278 18035 22330
rect 18059 22278 18073 22330
rect 18073 22278 18085 22330
rect 18085 22278 18115 22330
rect 18139 22278 18149 22330
rect 18149 22278 18195 22330
rect 17899 22276 17955 22278
rect 17979 22276 18035 22278
rect 18059 22276 18115 22278
rect 18139 22276 18195 22278
rect 17038 19780 17094 19816
rect 17038 19760 17040 19780
rect 17040 19760 17092 19780
rect 17092 19760 17094 19780
rect 16946 18808 17002 18864
rect 16394 10376 16450 10432
rect 16118 8492 16174 8528
rect 16118 8472 16120 8492
rect 16120 8472 16172 8492
rect 16172 8472 16174 8492
rect 15750 6740 15752 6760
rect 15752 6740 15804 6760
rect 15804 6740 15806 6760
rect 15750 6704 15806 6740
rect 15658 6568 15714 6624
rect 14510 2202 14566 2204
rect 14590 2202 14646 2204
rect 14670 2202 14726 2204
rect 14750 2202 14806 2204
rect 14510 2150 14556 2202
rect 14556 2150 14566 2202
rect 14590 2150 14620 2202
rect 14620 2150 14632 2202
rect 14632 2150 14646 2202
rect 14670 2150 14684 2202
rect 14684 2150 14696 2202
rect 14696 2150 14726 2202
rect 14750 2150 14760 2202
rect 14760 2150 14806 2202
rect 14510 2148 14566 2150
rect 14590 2148 14646 2150
rect 14670 2148 14726 2150
rect 14750 2148 14806 2150
rect 16210 7248 16266 7304
rect 16486 7248 16542 7304
rect 17314 16632 17370 16688
rect 17222 16496 17278 16552
rect 16854 13912 16910 13968
rect 17130 13368 17186 13424
rect 16670 10124 16726 10160
rect 16670 10104 16672 10124
rect 16672 10104 16724 10124
rect 16724 10104 16726 10124
rect 16578 6840 16634 6896
rect 17899 21242 17955 21244
rect 17979 21242 18035 21244
rect 18059 21242 18115 21244
rect 18139 21242 18195 21244
rect 17899 21190 17945 21242
rect 17945 21190 17955 21242
rect 17979 21190 18009 21242
rect 18009 21190 18021 21242
rect 18021 21190 18035 21242
rect 18059 21190 18073 21242
rect 18073 21190 18085 21242
rect 18085 21190 18115 21242
rect 18139 21190 18149 21242
rect 18149 21190 18195 21242
rect 17899 21188 17955 21190
rect 17979 21188 18035 21190
rect 18059 21188 18115 21190
rect 18139 21188 18195 21190
rect 17866 20848 17922 20904
rect 17899 20154 17955 20156
rect 17979 20154 18035 20156
rect 18059 20154 18115 20156
rect 18139 20154 18195 20156
rect 17899 20102 17945 20154
rect 17945 20102 17955 20154
rect 17979 20102 18009 20154
rect 18009 20102 18021 20154
rect 18021 20102 18035 20154
rect 18059 20102 18073 20154
rect 18073 20102 18085 20154
rect 18085 20102 18115 20154
rect 18139 20102 18149 20154
rect 18149 20102 18195 20154
rect 17899 20100 17955 20102
rect 17979 20100 18035 20102
rect 18059 20100 18115 20102
rect 18139 20100 18195 20102
rect 18694 23704 18750 23760
rect 18510 22072 18566 22128
rect 17899 19066 17955 19068
rect 17979 19066 18035 19068
rect 18059 19066 18115 19068
rect 18139 19066 18195 19068
rect 17899 19014 17945 19066
rect 17945 19014 17955 19066
rect 17979 19014 18009 19066
rect 18009 19014 18021 19066
rect 18021 19014 18035 19066
rect 18059 19014 18073 19066
rect 18073 19014 18085 19066
rect 18085 19014 18115 19066
rect 18139 19014 18149 19066
rect 18149 19014 18195 19066
rect 17899 19012 17955 19014
rect 17979 19012 18035 19014
rect 18059 19012 18115 19014
rect 18139 19012 18195 19014
rect 17498 17720 17554 17776
rect 17498 16632 17554 16688
rect 17899 17978 17955 17980
rect 17979 17978 18035 17980
rect 18059 17978 18115 17980
rect 18139 17978 18195 17980
rect 17899 17926 17945 17978
rect 17945 17926 17955 17978
rect 17979 17926 18009 17978
rect 18009 17926 18021 17978
rect 18021 17926 18035 17978
rect 18059 17926 18073 17978
rect 18073 17926 18085 17978
rect 18085 17926 18115 17978
rect 18139 17926 18149 17978
rect 18149 17926 18195 17978
rect 17899 17924 17955 17926
rect 17979 17924 18035 17926
rect 18059 17924 18115 17926
rect 18139 17924 18195 17926
rect 17682 17196 17738 17232
rect 17682 17176 17684 17196
rect 17684 17176 17736 17196
rect 17736 17176 17738 17196
rect 17774 17040 17830 17096
rect 17899 16890 17955 16892
rect 17979 16890 18035 16892
rect 18059 16890 18115 16892
rect 18139 16890 18195 16892
rect 17899 16838 17945 16890
rect 17945 16838 17955 16890
rect 17979 16838 18009 16890
rect 18009 16838 18021 16890
rect 18021 16838 18035 16890
rect 18059 16838 18073 16890
rect 18073 16838 18085 16890
rect 18085 16838 18115 16890
rect 18139 16838 18149 16890
rect 18149 16838 18195 16890
rect 17899 16836 17955 16838
rect 17979 16836 18035 16838
rect 18059 16836 18115 16838
rect 18139 16836 18195 16838
rect 17899 15802 17955 15804
rect 17979 15802 18035 15804
rect 18059 15802 18115 15804
rect 18139 15802 18195 15804
rect 17899 15750 17945 15802
rect 17945 15750 17955 15802
rect 17979 15750 18009 15802
rect 18009 15750 18021 15802
rect 18021 15750 18035 15802
rect 18059 15750 18073 15802
rect 18073 15750 18085 15802
rect 18085 15750 18115 15802
rect 18139 15750 18149 15802
rect 18149 15750 18195 15802
rect 17899 15748 17955 15750
rect 17979 15748 18035 15750
rect 18059 15748 18115 15750
rect 18139 15748 18195 15750
rect 17899 14714 17955 14716
rect 17979 14714 18035 14716
rect 18059 14714 18115 14716
rect 18139 14714 18195 14716
rect 17899 14662 17945 14714
rect 17945 14662 17955 14714
rect 17979 14662 18009 14714
rect 18009 14662 18021 14714
rect 18021 14662 18035 14714
rect 18059 14662 18073 14714
rect 18073 14662 18085 14714
rect 18085 14662 18115 14714
rect 18139 14662 18149 14714
rect 18149 14662 18195 14714
rect 17899 14660 17955 14662
rect 17979 14660 18035 14662
rect 18059 14660 18115 14662
rect 18139 14660 18195 14662
rect 17406 12688 17462 12744
rect 17406 12180 17408 12200
rect 17408 12180 17460 12200
rect 17460 12180 17462 12200
rect 17406 12144 17462 12180
rect 17314 11464 17370 11520
rect 17038 9560 17094 9616
rect 17222 10412 17224 10432
rect 17224 10412 17276 10432
rect 17276 10412 17278 10432
rect 17222 10376 17278 10412
rect 17130 7248 17186 7304
rect 17038 6704 17094 6760
rect 18142 13912 18198 13968
rect 18510 17584 18566 17640
rect 19246 22888 19302 22944
rect 19154 21256 19210 21312
rect 17899 13626 17955 13628
rect 17979 13626 18035 13628
rect 18059 13626 18115 13628
rect 18139 13626 18195 13628
rect 17899 13574 17945 13626
rect 17945 13574 17955 13626
rect 17979 13574 18009 13626
rect 18009 13574 18021 13626
rect 18021 13574 18035 13626
rect 18059 13574 18073 13626
rect 18073 13574 18085 13626
rect 18085 13574 18115 13626
rect 18139 13574 18149 13626
rect 18149 13574 18195 13626
rect 17899 13572 17955 13574
rect 17979 13572 18035 13574
rect 18059 13572 18115 13574
rect 18139 13572 18195 13574
rect 17899 12538 17955 12540
rect 17979 12538 18035 12540
rect 18059 12538 18115 12540
rect 18139 12538 18195 12540
rect 17899 12486 17945 12538
rect 17945 12486 17955 12538
rect 17979 12486 18009 12538
rect 18009 12486 18021 12538
rect 18021 12486 18035 12538
rect 18059 12486 18073 12538
rect 18073 12486 18085 12538
rect 18085 12486 18115 12538
rect 18139 12486 18149 12538
rect 18149 12486 18195 12538
rect 17899 12484 17955 12486
rect 17979 12484 18035 12486
rect 18059 12484 18115 12486
rect 18139 12484 18195 12486
rect 17682 12280 17738 12336
rect 17590 11600 17646 11656
rect 17314 6568 17370 6624
rect 17498 9424 17554 9480
rect 17899 11450 17955 11452
rect 17979 11450 18035 11452
rect 18059 11450 18115 11452
rect 18139 11450 18195 11452
rect 17899 11398 17945 11450
rect 17945 11398 17955 11450
rect 17979 11398 18009 11450
rect 18009 11398 18021 11450
rect 18021 11398 18035 11450
rect 18059 11398 18073 11450
rect 18073 11398 18085 11450
rect 18085 11398 18115 11450
rect 18139 11398 18149 11450
rect 18149 11398 18195 11450
rect 17899 11396 17955 11398
rect 17979 11396 18035 11398
rect 18059 11396 18115 11398
rect 18139 11396 18195 11398
rect 17498 7520 17554 7576
rect 17682 5616 17738 5672
rect 17498 5108 17500 5128
rect 17500 5108 17552 5128
rect 17552 5108 17554 5128
rect 17498 5072 17554 5108
rect 17899 10362 17955 10364
rect 17979 10362 18035 10364
rect 18059 10362 18115 10364
rect 18139 10362 18195 10364
rect 17899 10310 17945 10362
rect 17945 10310 17955 10362
rect 17979 10310 18009 10362
rect 18009 10310 18021 10362
rect 18021 10310 18035 10362
rect 18059 10310 18073 10362
rect 18073 10310 18085 10362
rect 18085 10310 18115 10362
rect 18139 10310 18149 10362
rect 18149 10310 18195 10362
rect 17899 10308 17955 10310
rect 17979 10308 18035 10310
rect 18059 10308 18115 10310
rect 18139 10308 18195 10310
rect 18602 13252 18658 13288
rect 18602 13232 18604 13252
rect 18604 13232 18656 13252
rect 18656 13232 18658 13252
rect 18510 13096 18566 13152
rect 18418 12144 18474 12200
rect 18694 10648 18750 10704
rect 17899 9274 17955 9276
rect 17979 9274 18035 9276
rect 18059 9274 18115 9276
rect 18139 9274 18195 9276
rect 17899 9222 17945 9274
rect 17945 9222 17955 9274
rect 17979 9222 18009 9274
rect 18009 9222 18021 9274
rect 18021 9222 18035 9274
rect 18059 9222 18073 9274
rect 18073 9222 18085 9274
rect 18085 9222 18115 9274
rect 18139 9222 18149 9274
rect 18149 9222 18195 9274
rect 17899 9220 17955 9222
rect 17979 9220 18035 9222
rect 18059 9220 18115 9222
rect 18139 9220 18195 9222
rect 18326 9424 18382 9480
rect 17899 8186 17955 8188
rect 17979 8186 18035 8188
rect 18059 8186 18115 8188
rect 18139 8186 18195 8188
rect 17899 8134 17945 8186
rect 17945 8134 17955 8186
rect 17979 8134 18009 8186
rect 18009 8134 18021 8186
rect 18021 8134 18035 8186
rect 18059 8134 18073 8186
rect 18073 8134 18085 8186
rect 18085 8134 18115 8186
rect 18139 8134 18149 8186
rect 18149 8134 18195 8186
rect 17899 8132 17955 8134
rect 17979 8132 18035 8134
rect 18059 8132 18115 8134
rect 18139 8132 18195 8134
rect 17958 7928 18014 7984
rect 18142 7520 18198 7576
rect 17899 7098 17955 7100
rect 17979 7098 18035 7100
rect 18059 7098 18115 7100
rect 18139 7098 18195 7100
rect 17899 7046 17945 7098
rect 17945 7046 17955 7098
rect 17979 7046 18009 7098
rect 18009 7046 18021 7098
rect 18021 7046 18035 7098
rect 18059 7046 18073 7098
rect 18073 7046 18085 7098
rect 18085 7046 18115 7098
rect 18139 7046 18149 7098
rect 18149 7046 18195 7098
rect 17899 7044 17955 7046
rect 17979 7044 18035 7046
rect 18059 7044 18115 7046
rect 18139 7044 18195 7046
rect 18602 9424 18658 9480
rect 18786 8472 18842 8528
rect 18326 6704 18382 6760
rect 17899 6010 17955 6012
rect 17979 6010 18035 6012
rect 18059 6010 18115 6012
rect 18139 6010 18195 6012
rect 17899 5958 17945 6010
rect 17945 5958 17955 6010
rect 17979 5958 18009 6010
rect 18009 5958 18021 6010
rect 18021 5958 18035 6010
rect 18059 5958 18073 6010
rect 18073 5958 18085 6010
rect 18085 5958 18115 6010
rect 18139 5958 18149 6010
rect 18149 5958 18195 6010
rect 17899 5956 17955 5958
rect 17979 5956 18035 5958
rect 18059 5956 18115 5958
rect 18139 5956 18195 5958
rect 17899 4922 17955 4924
rect 17979 4922 18035 4924
rect 18059 4922 18115 4924
rect 18139 4922 18195 4924
rect 17899 4870 17945 4922
rect 17945 4870 17955 4922
rect 17979 4870 18009 4922
rect 18009 4870 18021 4922
rect 18021 4870 18035 4922
rect 18059 4870 18073 4922
rect 18073 4870 18085 4922
rect 18085 4870 18115 4922
rect 18139 4870 18149 4922
rect 18149 4870 18195 4922
rect 17899 4868 17955 4870
rect 17979 4868 18035 4870
rect 18059 4868 18115 4870
rect 18139 4868 18195 4870
rect 17899 3834 17955 3836
rect 17979 3834 18035 3836
rect 18059 3834 18115 3836
rect 18139 3834 18195 3836
rect 17899 3782 17945 3834
rect 17945 3782 17955 3834
rect 17979 3782 18009 3834
rect 18009 3782 18021 3834
rect 18021 3782 18035 3834
rect 18059 3782 18073 3834
rect 18073 3782 18085 3834
rect 18085 3782 18115 3834
rect 18139 3782 18149 3834
rect 18149 3782 18195 3834
rect 17899 3780 17955 3782
rect 17979 3780 18035 3782
rect 18059 3780 18115 3782
rect 18139 3780 18195 3782
rect 17958 3576 18014 3632
rect 18142 3304 18198 3360
rect 19062 17720 19118 17776
rect 19246 16632 19302 16688
rect 19246 15816 19302 15872
rect 19246 14184 19302 14240
rect 20166 20712 20222 20768
rect 20626 20748 20628 20768
rect 20628 20748 20680 20768
rect 20680 20748 20682 20768
rect 20626 20712 20682 20748
rect 19706 19488 19762 19544
rect 19890 19352 19946 19408
rect 19246 11464 19302 11520
rect 19154 8492 19210 8528
rect 19154 8472 19156 8492
rect 19156 8472 19208 8492
rect 19208 8472 19210 8492
rect 19062 8336 19118 8392
rect 18786 6704 18842 6760
rect 17899 2746 17955 2748
rect 17979 2746 18035 2748
rect 18059 2746 18115 2748
rect 18139 2746 18195 2748
rect 17899 2694 17945 2746
rect 17945 2694 17955 2746
rect 17979 2694 18009 2746
rect 18009 2694 18021 2746
rect 18021 2694 18035 2746
rect 18059 2694 18073 2746
rect 18073 2694 18085 2746
rect 18085 2694 18115 2746
rect 18139 2694 18149 2746
rect 18149 2694 18195 2746
rect 17899 2692 17955 2694
rect 17979 2692 18035 2694
rect 18059 2692 18115 2694
rect 18139 2692 18195 2694
rect 17590 856 17646 912
rect 18878 6160 18934 6216
rect 18878 2488 18934 2544
rect 19890 15000 19946 15056
rect 20626 19660 20628 19680
rect 20628 19660 20680 19680
rect 20680 19660 20682 19680
rect 20626 19624 20682 19660
rect 20442 18536 20498 18592
rect 20718 12280 20774 12336
rect 20718 8744 20774 8800
rect 19246 6024 19302 6080
rect 19338 5752 19394 5808
rect 19522 3460 19578 3496
rect 19522 3440 19524 3460
rect 19524 3440 19576 3460
rect 19576 3440 19578 3460
rect 19982 5908 20038 5944
rect 19982 5888 19984 5908
rect 19984 5888 20036 5908
rect 20036 5888 20038 5908
rect 20534 7112 20590 7168
rect 20534 5208 20590 5264
rect 20718 4392 20774 4448
rect 20258 4140 20314 4176
rect 20258 4120 20260 4140
rect 20260 4120 20312 4140
rect 20312 4120 20314 4140
rect 19982 1672 20038 1728
rect 16946 40 17002 96
<< metal3 >>
rect 0 24578 800 24608
rect 3141 24578 3207 24581
rect 0 24576 3207 24578
rect 0 24520 3146 24576
rect 3202 24520 3207 24576
rect 0 24518 3207 24520
rect 0 24488 800 24518
rect 3141 24515 3207 24518
rect 0 23762 800 23792
rect 2773 23762 2839 23765
rect 0 23760 2839 23762
rect 0 23704 2778 23760
rect 2834 23704 2839 23760
rect 0 23702 2839 23704
rect 0 23672 800 23702
rect 2773 23699 2839 23702
rect 18689 23762 18755 23765
rect 21767 23762 22567 23792
rect 18689 23760 22567 23762
rect 18689 23704 18694 23760
rect 18750 23704 22567 23760
rect 18689 23702 22567 23704
rect 18689 23699 18755 23702
rect 21767 23672 22567 23702
rect 0 22946 800 22976
rect 2313 22946 2379 22949
rect 0 22944 2379 22946
rect 0 22888 2318 22944
rect 2374 22888 2379 22944
rect 0 22886 2379 22888
rect 0 22856 800 22886
rect 2313 22883 2379 22886
rect 19241 22946 19307 22949
rect 21767 22946 22567 22976
rect 19241 22944 22567 22946
rect 19241 22888 19246 22944
rect 19302 22888 22567 22944
rect 19241 22886 22567 22888
rect 19241 22883 19307 22886
rect 21767 22856 22567 22886
rect 4332 22336 4652 22337
rect 4332 22272 4340 22336
rect 4404 22272 4420 22336
rect 4484 22272 4500 22336
rect 4564 22272 4580 22336
rect 4644 22272 4652 22336
rect 4332 22271 4652 22272
rect 11110 22336 11430 22337
rect 11110 22272 11118 22336
rect 11182 22272 11198 22336
rect 11262 22272 11278 22336
rect 11342 22272 11358 22336
rect 11422 22272 11430 22336
rect 11110 22271 11430 22272
rect 17887 22336 18207 22337
rect 17887 22272 17895 22336
rect 17959 22272 17975 22336
rect 18039 22272 18055 22336
rect 18119 22272 18135 22336
rect 18199 22272 18207 22336
rect 17887 22271 18207 22272
rect 0 22130 800 22160
rect 1853 22130 1919 22133
rect 0 22128 1919 22130
rect 0 22072 1858 22128
rect 1914 22072 1919 22128
rect 0 22070 1919 22072
rect 0 22040 800 22070
rect 1853 22067 1919 22070
rect 18505 22130 18571 22133
rect 21767 22130 22567 22160
rect 18505 22128 22567 22130
rect 18505 22072 18510 22128
rect 18566 22072 22567 22128
rect 18505 22070 22567 22072
rect 18505 22067 18571 22070
rect 21767 22040 22567 22070
rect 7721 21792 8041 21793
rect 7721 21728 7729 21792
rect 7793 21728 7809 21792
rect 7873 21728 7889 21792
rect 7953 21728 7969 21792
rect 8033 21728 8041 21792
rect 7721 21727 8041 21728
rect 14498 21792 14818 21793
rect 14498 21728 14506 21792
rect 14570 21728 14586 21792
rect 14650 21728 14666 21792
rect 14730 21728 14746 21792
rect 14810 21728 14818 21792
rect 14498 21727 14818 21728
rect 10041 21450 10107 21453
rect 14365 21450 14431 21453
rect 10041 21448 14431 21450
rect 10041 21392 10046 21448
rect 10102 21392 14370 21448
rect 14426 21392 14431 21448
rect 10041 21390 14431 21392
rect 10041 21387 10107 21390
rect 14365 21387 14431 21390
rect 19149 21314 19215 21317
rect 21767 21314 22567 21344
rect 19149 21312 22567 21314
rect 19149 21256 19154 21312
rect 19210 21256 22567 21312
rect 19149 21254 22567 21256
rect 19149 21251 19215 21254
rect 4332 21248 4652 21249
rect 4332 21184 4340 21248
rect 4404 21184 4420 21248
rect 4484 21184 4500 21248
rect 4564 21184 4580 21248
rect 4644 21184 4652 21248
rect 4332 21183 4652 21184
rect 11110 21248 11430 21249
rect 11110 21184 11118 21248
rect 11182 21184 11198 21248
rect 11262 21184 11278 21248
rect 11342 21184 11358 21248
rect 11422 21184 11430 21248
rect 11110 21183 11430 21184
rect 17887 21248 18207 21249
rect 17887 21184 17895 21248
rect 17959 21184 17975 21248
rect 18039 21184 18055 21248
rect 18119 21184 18135 21248
rect 18199 21184 18207 21248
rect 21767 21224 22567 21254
rect 17887 21183 18207 21184
rect 0 21042 800 21072
rect 3233 21042 3299 21045
rect 0 21040 3299 21042
rect 0 20984 3238 21040
rect 3294 20984 3299 21040
rect 0 20982 3299 20984
rect 0 20952 800 20982
rect 3233 20979 3299 20982
rect 10133 21042 10199 21045
rect 11053 21042 11119 21045
rect 10133 21040 11119 21042
rect 10133 20984 10138 21040
rect 10194 20984 11058 21040
rect 11114 20984 11119 21040
rect 10133 20982 11119 20984
rect 10133 20979 10199 20982
rect 11053 20979 11119 20982
rect 12065 21042 12131 21045
rect 16481 21042 16547 21045
rect 16757 21042 16823 21045
rect 12065 21040 16823 21042
rect 12065 20984 12070 21040
rect 12126 20984 16486 21040
rect 16542 20984 16762 21040
rect 16818 20984 16823 21040
rect 12065 20982 16823 20984
rect 12065 20979 12131 20982
rect 16481 20979 16547 20982
rect 16757 20979 16823 20982
rect 10777 20906 10843 20909
rect 17861 20906 17927 20909
rect 10777 20904 17927 20906
rect 10777 20848 10782 20904
rect 10838 20848 17866 20904
rect 17922 20848 17927 20904
rect 10777 20846 17927 20848
rect 10777 20843 10843 20846
rect 17861 20843 17927 20846
rect 10041 20770 10107 20773
rect 12065 20770 12131 20773
rect 10041 20768 12131 20770
rect 10041 20712 10046 20768
rect 10102 20712 12070 20768
rect 12126 20712 12131 20768
rect 10041 20710 12131 20712
rect 10041 20707 10107 20710
rect 12065 20707 12131 20710
rect 20161 20770 20227 20773
rect 20294 20770 20300 20772
rect 20161 20768 20300 20770
rect 20161 20712 20166 20768
rect 20222 20712 20300 20768
rect 20161 20710 20300 20712
rect 20161 20707 20227 20710
rect 20294 20708 20300 20710
rect 20364 20708 20370 20772
rect 20478 20708 20484 20772
rect 20548 20770 20554 20772
rect 20621 20770 20687 20773
rect 20548 20768 20687 20770
rect 20548 20712 20626 20768
rect 20682 20712 20687 20768
rect 20548 20710 20687 20712
rect 20548 20708 20554 20710
rect 20621 20707 20687 20710
rect 7721 20704 8041 20705
rect 7721 20640 7729 20704
rect 7793 20640 7809 20704
rect 7873 20640 7889 20704
rect 7953 20640 7969 20704
rect 8033 20640 8041 20704
rect 7721 20639 8041 20640
rect 14498 20704 14818 20705
rect 14498 20640 14506 20704
rect 14570 20640 14586 20704
rect 14650 20640 14666 20704
rect 14730 20640 14746 20704
rect 14810 20640 14818 20704
rect 14498 20639 14818 20640
rect 5809 20634 5875 20637
rect 7373 20634 7439 20637
rect 5809 20632 7439 20634
rect 5809 20576 5814 20632
rect 5870 20576 7378 20632
rect 7434 20576 7439 20632
rect 5809 20574 7439 20576
rect 5809 20571 5875 20574
rect 7373 20571 7439 20574
rect 5349 20498 5415 20501
rect 6269 20498 6335 20501
rect 5349 20496 6335 20498
rect 5349 20440 5354 20496
rect 5410 20440 6274 20496
rect 6330 20440 6335 20496
rect 5349 20438 6335 20440
rect 5349 20435 5415 20438
rect 6269 20435 6335 20438
rect 6637 20498 6703 20501
rect 8753 20498 8819 20501
rect 6637 20496 8819 20498
rect 6637 20440 6642 20496
rect 6698 20440 8758 20496
rect 8814 20440 8819 20496
rect 6637 20438 8819 20440
rect 6637 20435 6703 20438
rect 8753 20435 8819 20438
rect 5349 20362 5415 20365
rect 6085 20362 6151 20365
rect 5349 20360 6151 20362
rect 5349 20304 5354 20360
rect 5410 20304 6090 20360
rect 6146 20304 6151 20360
rect 5349 20302 6151 20304
rect 5349 20299 5415 20302
rect 6085 20299 6151 20302
rect 0 20226 800 20256
rect 1577 20226 1643 20229
rect 0 20224 1643 20226
rect 0 20168 1582 20224
rect 1638 20168 1643 20224
rect 0 20166 1643 20168
rect 0 20136 800 20166
rect 1577 20163 1643 20166
rect 4332 20160 4652 20161
rect 4332 20096 4340 20160
rect 4404 20096 4420 20160
rect 4484 20096 4500 20160
rect 4564 20096 4580 20160
rect 4644 20096 4652 20160
rect 4332 20095 4652 20096
rect 11110 20160 11430 20161
rect 11110 20096 11118 20160
rect 11182 20096 11198 20160
rect 11262 20096 11278 20160
rect 11342 20096 11358 20160
rect 11422 20096 11430 20160
rect 11110 20095 11430 20096
rect 17887 20160 18207 20161
rect 17887 20096 17895 20160
rect 17959 20096 17975 20160
rect 18039 20096 18055 20160
rect 18119 20096 18135 20160
rect 18199 20096 18207 20160
rect 21767 20136 22567 20256
rect 17887 20095 18207 20096
rect 11513 20090 11579 20093
rect 12893 20090 12959 20093
rect 11513 20088 12959 20090
rect 11513 20032 11518 20088
rect 11574 20032 12898 20088
rect 12954 20032 12959 20088
rect 11513 20030 12959 20032
rect 11513 20027 11579 20030
rect 12893 20027 12959 20030
rect 7557 19818 7623 19821
rect 17033 19818 17099 19821
rect 7557 19816 17099 19818
rect 7557 19760 7562 19816
rect 7618 19760 17038 19816
rect 17094 19760 17099 19816
rect 7557 19758 17099 19760
rect 7557 19755 7623 19758
rect 17033 19755 17099 19758
rect 19926 19620 19932 19684
rect 19996 19682 20002 19684
rect 20621 19682 20687 19685
rect 19996 19680 20687 19682
rect 19996 19624 20626 19680
rect 20682 19624 20687 19680
rect 19996 19622 20687 19624
rect 19996 19620 20002 19622
rect 20621 19619 20687 19622
rect 7721 19616 8041 19617
rect 7721 19552 7729 19616
rect 7793 19552 7809 19616
rect 7873 19552 7889 19616
rect 7953 19552 7969 19616
rect 8033 19552 8041 19616
rect 7721 19551 8041 19552
rect 14498 19616 14818 19617
rect 14498 19552 14506 19616
rect 14570 19552 14586 19616
rect 14650 19552 14666 19616
rect 14730 19552 14746 19616
rect 14810 19552 14818 19616
rect 14498 19551 14818 19552
rect 9765 19546 9831 19549
rect 12341 19546 12407 19549
rect 13721 19546 13787 19549
rect 9765 19544 12082 19546
rect 9765 19488 9770 19544
rect 9826 19488 12082 19544
rect 9765 19486 12082 19488
rect 9765 19483 9831 19486
rect 0 19410 800 19440
rect 1393 19410 1459 19413
rect 0 19408 1459 19410
rect 0 19352 1398 19408
rect 1454 19352 1459 19408
rect 0 19350 1459 19352
rect 0 19320 800 19350
rect 1393 19347 1459 19350
rect 2313 19410 2379 19413
rect 4797 19410 4863 19413
rect 2313 19408 4863 19410
rect 2313 19352 2318 19408
rect 2374 19352 4802 19408
rect 4858 19352 4863 19408
rect 2313 19350 4863 19352
rect 2313 19347 2379 19350
rect 4797 19347 4863 19350
rect 9305 19410 9371 19413
rect 11881 19410 11947 19413
rect 9305 19408 11947 19410
rect 9305 19352 9310 19408
rect 9366 19352 11886 19408
rect 11942 19352 11947 19408
rect 9305 19350 11947 19352
rect 12022 19410 12082 19486
rect 12341 19544 13787 19546
rect 12341 19488 12346 19544
rect 12402 19488 13726 19544
rect 13782 19488 13787 19544
rect 12341 19486 13787 19488
rect 12341 19483 12407 19486
rect 13721 19483 13787 19486
rect 19701 19546 19767 19549
rect 20110 19546 20116 19548
rect 19701 19544 20116 19546
rect 19701 19488 19706 19544
rect 19762 19488 20116 19544
rect 19701 19486 20116 19488
rect 19701 19483 19767 19486
rect 20110 19484 20116 19486
rect 20180 19484 20186 19548
rect 12801 19410 12867 19413
rect 12022 19408 12867 19410
rect 12022 19352 12806 19408
rect 12862 19352 12867 19408
rect 12022 19350 12867 19352
rect 9305 19347 9371 19350
rect 11881 19347 11947 19350
rect 12801 19347 12867 19350
rect 19885 19410 19951 19413
rect 21767 19410 22567 19440
rect 19885 19408 22567 19410
rect 19885 19352 19890 19408
rect 19946 19352 22567 19408
rect 19885 19350 22567 19352
rect 19885 19347 19951 19350
rect 21767 19320 22567 19350
rect 3877 19274 3943 19277
rect 4245 19274 4311 19277
rect 3877 19272 4311 19274
rect 3877 19216 3882 19272
rect 3938 19216 4250 19272
rect 4306 19216 4311 19272
rect 3877 19214 4311 19216
rect 3877 19211 3943 19214
rect 4245 19211 4311 19214
rect 14917 19276 14983 19277
rect 14917 19272 14964 19276
rect 15028 19274 15034 19276
rect 14917 19216 14922 19272
rect 14917 19212 14964 19216
rect 15028 19214 15074 19274
rect 15028 19212 15034 19214
rect 14917 19211 14983 19212
rect 4332 19072 4652 19073
rect 4332 19008 4340 19072
rect 4404 19008 4420 19072
rect 4484 19008 4500 19072
rect 4564 19008 4580 19072
rect 4644 19008 4652 19072
rect 4332 19007 4652 19008
rect 11110 19072 11430 19073
rect 11110 19008 11118 19072
rect 11182 19008 11198 19072
rect 11262 19008 11278 19072
rect 11342 19008 11358 19072
rect 11422 19008 11430 19072
rect 11110 19007 11430 19008
rect 17887 19072 18207 19073
rect 17887 19008 17895 19072
rect 17959 19008 17975 19072
rect 18039 19008 18055 19072
rect 18119 19008 18135 19072
rect 18199 19008 18207 19072
rect 17887 19007 18207 19008
rect 10777 18866 10843 18869
rect 12525 18866 12591 18869
rect 13169 18866 13235 18869
rect 16941 18866 17007 18869
rect 10777 18864 17007 18866
rect 10777 18808 10782 18864
rect 10838 18808 12530 18864
rect 12586 18808 13174 18864
rect 13230 18808 16946 18864
rect 17002 18808 17007 18864
rect 10777 18806 17007 18808
rect 10777 18803 10843 18806
rect 12525 18803 12591 18806
rect 13169 18803 13235 18806
rect 16941 18803 17007 18806
rect 6729 18730 6795 18733
rect 7189 18730 7255 18733
rect 6729 18728 7255 18730
rect 6729 18672 6734 18728
rect 6790 18672 7194 18728
rect 7250 18672 7255 18728
rect 6729 18670 7255 18672
rect 6729 18667 6795 18670
rect 7189 18667 7255 18670
rect 0 18594 800 18624
rect 1669 18594 1735 18597
rect 0 18592 1735 18594
rect 0 18536 1674 18592
rect 1730 18536 1735 18592
rect 0 18534 1735 18536
rect 0 18504 800 18534
rect 1669 18531 1735 18534
rect 20437 18594 20503 18597
rect 21767 18594 22567 18624
rect 20437 18592 22567 18594
rect 20437 18536 20442 18592
rect 20498 18536 22567 18592
rect 20437 18534 22567 18536
rect 20437 18531 20503 18534
rect 7721 18528 8041 18529
rect 7721 18464 7729 18528
rect 7793 18464 7809 18528
rect 7873 18464 7889 18528
rect 7953 18464 7969 18528
rect 8033 18464 8041 18528
rect 7721 18463 8041 18464
rect 14498 18528 14818 18529
rect 14498 18464 14506 18528
rect 14570 18464 14586 18528
rect 14650 18464 14666 18528
rect 14730 18464 14746 18528
rect 14810 18464 14818 18528
rect 21767 18504 22567 18534
rect 14498 18463 14818 18464
rect 11881 18322 11947 18325
rect 16573 18322 16639 18325
rect 11881 18320 16639 18322
rect 11881 18264 11886 18320
rect 11942 18264 16578 18320
rect 16634 18264 16639 18320
rect 11881 18262 16639 18264
rect 11881 18259 11947 18262
rect 16573 18259 16639 18262
rect 4332 17984 4652 17985
rect 4332 17920 4340 17984
rect 4404 17920 4420 17984
rect 4484 17920 4500 17984
rect 4564 17920 4580 17984
rect 4644 17920 4652 17984
rect 4332 17919 4652 17920
rect 11110 17984 11430 17985
rect 11110 17920 11118 17984
rect 11182 17920 11198 17984
rect 11262 17920 11278 17984
rect 11342 17920 11358 17984
rect 11422 17920 11430 17984
rect 11110 17919 11430 17920
rect 17887 17984 18207 17985
rect 17887 17920 17895 17984
rect 17959 17920 17975 17984
rect 18039 17920 18055 17984
rect 18119 17920 18135 17984
rect 18199 17920 18207 17984
rect 17887 17919 18207 17920
rect 12341 17914 12407 17917
rect 15469 17914 15535 17917
rect 12341 17912 15535 17914
rect 12341 17856 12346 17912
rect 12402 17856 15474 17912
rect 15530 17856 15535 17912
rect 12341 17854 15535 17856
rect 12341 17851 12407 17854
rect 15469 17851 15535 17854
rect 10225 17778 10291 17781
rect 17493 17778 17559 17781
rect 10225 17776 17559 17778
rect 10225 17720 10230 17776
rect 10286 17720 17498 17776
rect 17554 17720 17559 17776
rect 10225 17718 17559 17720
rect 10225 17715 10291 17718
rect 17493 17715 17559 17718
rect 19057 17778 19123 17781
rect 21767 17778 22567 17808
rect 19057 17776 22567 17778
rect 19057 17720 19062 17776
rect 19118 17720 22567 17776
rect 19057 17718 22567 17720
rect 19057 17715 19123 17718
rect 21767 17688 22567 17718
rect 4061 17642 4127 17645
rect 8477 17642 8543 17645
rect 4061 17640 8543 17642
rect 4061 17584 4066 17640
rect 4122 17584 8482 17640
rect 8538 17584 8543 17640
rect 4061 17582 8543 17584
rect 4061 17579 4127 17582
rect 8477 17579 8543 17582
rect 11513 17642 11579 17645
rect 18505 17642 18571 17645
rect 11513 17640 18571 17642
rect 11513 17584 11518 17640
rect 11574 17584 18510 17640
rect 18566 17584 18571 17640
rect 11513 17582 18571 17584
rect 11513 17579 11579 17582
rect 18505 17579 18571 17582
rect 0 17506 800 17536
rect 1853 17506 1919 17509
rect 0 17504 1919 17506
rect 0 17448 1858 17504
rect 1914 17448 1919 17504
rect 0 17446 1919 17448
rect 0 17416 800 17446
rect 1853 17443 1919 17446
rect 7721 17440 8041 17441
rect 7721 17376 7729 17440
rect 7793 17376 7809 17440
rect 7873 17376 7889 17440
rect 7953 17376 7969 17440
rect 8033 17376 8041 17440
rect 7721 17375 8041 17376
rect 14498 17440 14818 17441
rect 14498 17376 14506 17440
rect 14570 17376 14586 17440
rect 14650 17376 14666 17440
rect 14730 17376 14746 17440
rect 14810 17376 14818 17440
rect 14498 17375 14818 17376
rect 11973 17370 12039 17373
rect 13537 17370 13603 17373
rect 11973 17368 13603 17370
rect 11973 17312 11978 17368
rect 12034 17312 13542 17368
rect 13598 17312 13603 17368
rect 11973 17310 13603 17312
rect 11973 17307 12039 17310
rect 13537 17307 13603 17310
rect 3325 17234 3391 17237
rect 8845 17234 8911 17237
rect 3325 17232 8911 17234
rect 3325 17176 3330 17232
rect 3386 17176 8850 17232
rect 8906 17176 8911 17232
rect 3325 17174 8911 17176
rect 3325 17171 3391 17174
rect 8845 17171 8911 17174
rect 10777 17234 10843 17237
rect 17677 17234 17743 17237
rect 10777 17232 17743 17234
rect 10777 17176 10782 17232
rect 10838 17176 17682 17232
rect 17738 17176 17743 17232
rect 10777 17174 17743 17176
rect 10777 17171 10843 17174
rect 17677 17171 17743 17174
rect 12341 17098 12407 17101
rect 12801 17098 12867 17101
rect 12341 17096 12867 17098
rect 12341 17040 12346 17096
rect 12402 17040 12806 17096
rect 12862 17040 12867 17096
rect 12341 17038 12867 17040
rect 12341 17035 12407 17038
rect 12801 17035 12867 17038
rect 13721 17098 13787 17101
rect 17769 17098 17835 17101
rect 13721 17096 17835 17098
rect 13721 17040 13726 17096
rect 13782 17040 17774 17096
rect 17830 17040 17835 17096
rect 13721 17038 17835 17040
rect 13721 17035 13787 17038
rect 17769 17035 17835 17038
rect 4332 16896 4652 16897
rect 4332 16832 4340 16896
rect 4404 16832 4420 16896
rect 4484 16832 4500 16896
rect 4564 16832 4580 16896
rect 4644 16832 4652 16896
rect 4332 16831 4652 16832
rect 11110 16896 11430 16897
rect 11110 16832 11118 16896
rect 11182 16832 11198 16896
rect 11262 16832 11278 16896
rect 11342 16832 11358 16896
rect 11422 16832 11430 16896
rect 11110 16831 11430 16832
rect 17887 16896 18207 16897
rect 17887 16832 17895 16896
rect 17959 16832 17975 16896
rect 18039 16832 18055 16896
rect 18119 16832 18135 16896
rect 18199 16832 18207 16896
rect 17887 16831 18207 16832
rect 14181 16826 14247 16829
rect 14825 16826 14891 16829
rect 14181 16824 14891 16826
rect 14181 16768 14186 16824
rect 14242 16768 14830 16824
rect 14886 16768 14891 16824
rect 14181 16766 14891 16768
rect 14181 16763 14247 16766
rect 14825 16763 14891 16766
rect 0 16690 800 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 800 16630
rect 4061 16627 4127 16630
rect 10225 16690 10291 16693
rect 16573 16690 16639 16693
rect 17309 16690 17375 16693
rect 10225 16688 17375 16690
rect 10225 16632 10230 16688
rect 10286 16632 16578 16688
rect 16634 16632 17314 16688
rect 17370 16632 17375 16688
rect 10225 16630 17375 16632
rect 10225 16627 10291 16630
rect 16573 16627 16639 16630
rect 17309 16627 17375 16630
rect 17493 16690 17559 16693
rect 17718 16690 17724 16692
rect 17493 16688 17724 16690
rect 17493 16632 17498 16688
rect 17554 16632 17724 16688
rect 17493 16630 17724 16632
rect 17493 16627 17559 16630
rect 17718 16628 17724 16630
rect 17788 16628 17794 16692
rect 19241 16690 19307 16693
rect 21767 16690 22567 16720
rect 19241 16688 22567 16690
rect 19241 16632 19246 16688
rect 19302 16632 22567 16688
rect 19241 16630 22567 16632
rect 19241 16627 19307 16630
rect 21767 16600 22567 16630
rect 7281 16554 7347 16557
rect 9305 16556 9371 16557
rect 8150 16554 8156 16556
rect 7281 16552 8156 16554
rect 7281 16496 7286 16552
rect 7342 16496 8156 16552
rect 7281 16494 8156 16496
rect 7281 16491 7347 16494
rect 8150 16492 8156 16494
rect 8220 16492 8226 16556
rect 9254 16492 9260 16556
rect 9324 16554 9371 16556
rect 11973 16554 12039 16557
rect 17217 16554 17283 16557
rect 9324 16552 9416 16554
rect 9366 16496 9416 16552
rect 9324 16494 9416 16496
rect 11973 16552 17283 16554
rect 11973 16496 11978 16552
rect 12034 16496 17222 16552
rect 17278 16496 17283 16552
rect 11973 16494 17283 16496
rect 9324 16492 9371 16494
rect 9305 16491 9371 16492
rect 11973 16491 12039 16494
rect 17217 16491 17283 16494
rect 7721 16352 8041 16353
rect 7721 16288 7729 16352
rect 7793 16288 7809 16352
rect 7873 16288 7889 16352
rect 7953 16288 7969 16352
rect 8033 16288 8041 16352
rect 7721 16287 8041 16288
rect 14498 16352 14818 16353
rect 14498 16288 14506 16352
rect 14570 16288 14586 16352
rect 14650 16288 14666 16352
rect 14730 16288 14746 16352
rect 14810 16288 14818 16352
rect 14498 16287 14818 16288
rect 2681 16010 2747 16013
rect 6545 16010 6611 16013
rect 2681 16008 6611 16010
rect 2681 15952 2686 16008
rect 2742 15952 6550 16008
rect 6606 15952 6611 16008
rect 2681 15950 6611 15952
rect 2681 15947 2747 15950
rect 6545 15947 6611 15950
rect 10225 16010 10291 16013
rect 15745 16010 15811 16013
rect 10225 16008 15811 16010
rect 10225 15952 10230 16008
rect 10286 15952 15750 16008
rect 15806 15952 15811 16008
rect 10225 15950 15811 15952
rect 10225 15947 10291 15950
rect 15745 15947 15811 15950
rect 0 15874 800 15904
rect 2773 15874 2839 15877
rect 0 15872 2839 15874
rect 0 15816 2778 15872
rect 2834 15816 2839 15872
rect 0 15814 2839 15816
rect 0 15784 800 15814
rect 2773 15811 2839 15814
rect 19241 15874 19307 15877
rect 21767 15874 22567 15904
rect 19241 15872 22567 15874
rect 19241 15816 19246 15872
rect 19302 15816 22567 15872
rect 19241 15814 22567 15816
rect 19241 15811 19307 15814
rect 4332 15808 4652 15809
rect 4332 15744 4340 15808
rect 4404 15744 4420 15808
rect 4484 15744 4500 15808
rect 4564 15744 4580 15808
rect 4644 15744 4652 15808
rect 4332 15743 4652 15744
rect 11110 15808 11430 15809
rect 11110 15744 11118 15808
rect 11182 15744 11198 15808
rect 11262 15744 11278 15808
rect 11342 15744 11358 15808
rect 11422 15744 11430 15808
rect 11110 15743 11430 15744
rect 17887 15808 18207 15809
rect 17887 15744 17895 15808
rect 17959 15744 17975 15808
rect 18039 15744 18055 15808
rect 18119 15744 18135 15808
rect 18199 15744 18207 15808
rect 21767 15784 22567 15814
rect 17887 15743 18207 15744
rect 7721 15264 8041 15265
rect 7721 15200 7729 15264
rect 7793 15200 7809 15264
rect 7873 15200 7889 15264
rect 7953 15200 7969 15264
rect 8033 15200 8041 15264
rect 7721 15199 8041 15200
rect 14498 15264 14818 15265
rect 14498 15200 14506 15264
rect 14570 15200 14586 15264
rect 14650 15200 14666 15264
rect 14730 15200 14746 15264
rect 14810 15200 14818 15264
rect 14498 15199 14818 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 2773 15058 2839 15061
rect 3509 15058 3575 15061
rect 7741 15058 7807 15061
rect 16389 15058 16455 15061
rect 2773 15056 7807 15058
rect 2773 15000 2778 15056
rect 2834 15000 3514 15056
rect 3570 15000 7746 15056
rect 7802 15000 7807 15056
rect 2773 14998 7807 15000
rect 2773 14995 2839 14998
rect 3509 14995 3575 14998
rect 7741 14995 7807 14998
rect 16254 15056 16455 15058
rect 16254 15000 16394 15056
rect 16450 15000 16455 15056
rect 16254 14998 16455 15000
rect 9305 14922 9371 14925
rect 10685 14922 10751 14925
rect 9305 14920 10751 14922
rect 9305 14864 9310 14920
rect 9366 14864 10690 14920
rect 10746 14864 10751 14920
rect 9305 14862 10751 14864
rect 9305 14859 9371 14862
rect 10685 14859 10751 14862
rect 16113 14922 16179 14925
rect 16254 14922 16314 14998
rect 16389 14995 16455 14998
rect 19885 15058 19951 15061
rect 21767 15058 22567 15088
rect 19885 15056 22567 15058
rect 19885 15000 19890 15056
rect 19946 15000 22567 15056
rect 19885 14998 22567 15000
rect 19885 14995 19951 14998
rect 21767 14968 22567 14998
rect 16113 14920 16314 14922
rect 16113 14864 16118 14920
rect 16174 14864 16314 14920
rect 16113 14862 16314 14864
rect 16113 14859 16179 14862
rect 5717 14786 5783 14789
rect 6177 14786 6243 14789
rect 10961 14786 11027 14789
rect 5717 14784 11027 14786
rect 5717 14728 5722 14784
rect 5778 14728 6182 14784
rect 6238 14728 10966 14784
rect 11022 14728 11027 14784
rect 5717 14726 11027 14728
rect 5717 14723 5783 14726
rect 6177 14723 6243 14726
rect 10961 14723 11027 14726
rect 4332 14720 4652 14721
rect 4332 14656 4340 14720
rect 4404 14656 4420 14720
rect 4484 14656 4500 14720
rect 4564 14656 4580 14720
rect 4644 14656 4652 14720
rect 4332 14655 4652 14656
rect 11110 14720 11430 14721
rect 11110 14656 11118 14720
rect 11182 14656 11198 14720
rect 11262 14656 11278 14720
rect 11342 14656 11358 14720
rect 11422 14656 11430 14720
rect 11110 14655 11430 14656
rect 17887 14720 18207 14721
rect 17887 14656 17895 14720
rect 17959 14656 17975 14720
rect 18039 14656 18055 14720
rect 18119 14656 18135 14720
rect 18199 14656 18207 14720
rect 17887 14655 18207 14656
rect 9489 14650 9555 14653
rect 9446 14648 9555 14650
rect 9446 14592 9494 14648
rect 9550 14592 9555 14648
rect 9446 14587 9555 14592
rect 7721 14176 8041 14177
rect 7721 14112 7729 14176
rect 7793 14112 7809 14176
rect 7873 14112 7889 14176
rect 7953 14112 7969 14176
rect 8033 14112 8041 14176
rect 7721 14111 8041 14112
rect 9446 14109 9506 14587
rect 9673 14514 9739 14517
rect 10593 14514 10659 14517
rect 14733 14514 14799 14517
rect 9673 14512 14799 14514
rect 9673 14456 9678 14512
rect 9734 14456 10598 14512
rect 10654 14456 14738 14512
rect 14794 14456 14799 14512
rect 9673 14454 14799 14456
rect 9673 14451 9739 14454
rect 10593 14451 10659 14454
rect 14733 14451 14799 14454
rect 19241 14242 19307 14245
rect 21767 14242 22567 14272
rect 19241 14240 22567 14242
rect 19241 14184 19246 14240
rect 19302 14184 22567 14240
rect 19241 14182 22567 14184
rect 19241 14179 19307 14182
rect 14498 14176 14818 14177
rect 14498 14112 14506 14176
rect 14570 14112 14586 14176
rect 14650 14112 14666 14176
rect 14730 14112 14746 14176
rect 14810 14112 14818 14176
rect 21767 14152 22567 14182
rect 14498 14111 14818 14112
rect 5809 14106 5875 14109
rect 7465 14106 7531 14109
rect 9213 14108 9279 14109
rect 9213 14106 9260 14108
rect 5809 14104 7531 14106
rect 5809 14048 5814 14104
rect 5870 14048 7470 14104
rect 7526 14048 7531 14104
rect 5809 14046 7531 14048
rect 9168 14104 9260 14106
rect 9168 14048 9218 14104
rect 9168 14046 9260 14048
rect 5809 14043 5875 14046
rect 7465 14043 7531 14046
rect 9213 14044 9260 14046
rect 9324 14044 9330 14108
rect 9446 14104 9555 14109
rect 9446 14048 9494 14104
rect 9550 14048 9555 14104
rect 9446 14046 9555 14048
rect 9213 14043 9279 14044
rect 9489 14043 9555 14046
rect 0 13970 800 14000
rect 1669 13970 1735 13973
rect 0 13968 1735 13970
rect 0 13912 1674 13968
rect 1730 13912 1735 13968
rect 0 13910 1735 13912
rect 0 13880 800 13910
rect 1669 13907 1735 13910
rect 9949 13970 10015 13973
rect 16849 13970 16915 13973
rect 9949 13968 16915 13970
rect 9949 13912 9954 13968
rect 10010 13912 16854 13968
rect 16910 13912 16915 13968
rect 9949 13910 16915 13912
rect 9949 13907 10015 13910
rect 16849 13907 16915 13910
rect 17718 13908 17724 13972
rect 17788 13970 17794 13972
rect 18137 13970 18203 13973
rect 17788 13968 18203 13970
rect 17788 13912 18142 13968
rect 18198 13912 18203 13968
rect 17788 13910 18203 13912
rect 17788 13908 17794 13910
rect 15745 13834 15811 13837
rect 17726 13834 17786 13908
rect 18137 13907 18203 13910
rect 15745 13832 17786 13834
rect 15745 13776 15750 13832
rect 15806 13776 17786 13832
rect 15745 13774 17786 13776
rect 15745 13771 15811 13774
rect 4332 13632 4652 13633
rect 4332 13568 4340 13632
rect 4404 13568 4420 13632
rect 4484 13568 4500 13632
rect 4564 13568 4580 13632
rect 4644 13568 4652 13632
rect 4332 13567 4652 13568
rect 11110 13632 11430 13633
rect 11110 13568 11118 13632
rect 11182 13568 11198 13632
rect 11262 13568 11278 13632
rect 11342 13568 11358 13632
rect 11422 13568 11430 13632
rect 11110 13567 11430 13568
rect 17887 13632 18207 13633
rect 17887 13568 17895 13632
rect 17959 13568 17975 13632
rect 18039 13568 18055 13632
rect 18119 13568 18135 13632
rect 18199 13568 18207 13632
rect 17887 13567 18207 13568
rect 10133 13426 10199 13429
rect 12617 13426 12683 13429
rect 10133 13424 12683 13426
rect 10133 13368 10138 13424
rect 10194 13368 12622 13424
rect 12678 13368 12683 13424
rect 10133 13366 12683 13368
rect 10133 13363 10199 13366
rect 12617 13363 12683 13366
rect 14958 13364 14964 13428
rect 15028 13426 15034 13428
rect 15101 13426 15167 13429
rect 17125 13426 17191 13429
rect 15028 13424 17191 13426
rect 15028 13368 15106 13424
rect 15162 13368 17130 13424
rect 17186 13368 17191 13424
rect 15028 13366 17191 13368
rect 15028 13364 15034 13366
rect 15101 13363 15167 13366
rect 17125 13363 17191 13366
rect 15469 13290 15535 13293
rect 15653 13290 15719 13293
rect 18597 13290 18663 13293
rect 15469 13288 18663 13290
rect 15469 13232 15474 13288
rect 15530 13232 15658 13288
rect 15714 13232 18602 13288
rect 18658 13232 18663 13288
rect 15469 13230 18663 13232
rect 15469 13227 15535 13230
rect 15653 13227 15719 13230
rect 18597 13227 18663 13230
rect 0 13154 800 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 800 13094
rect 1577 13091 1643 13094
rect 18505 13154 18571 13157
rect 21767 13154 22567 13184
rect 18505 13152 22567 13154
rect 18505 13096 18510 13152
rect 18566 13096 22567 13152
rect 18505 13094 22567 13096
rect 18505 13091 18571 13094
rect 7721 13088 8041 13089
rect 7721 13024 7729 13088
rect 7793 13024 7809 13088
rect 7873 13024 7889 13088
rect 7953 13024 7969 13088
rect 8033 13024 8041 13088
rect 7721 13023 8041 13024
rect 14498 13088 14818 13089
rect 14498 13024 14506 13088
rect 14570 13024 14586 13088
rect 14650 13024 14666 13088
rect 14730 13024 14746 13088
rect 14810 13024 14818 13088
rect 21767 13064 22567 13094
rect 14498 13023 14818 13024
rect 8845 13018 8911 13021
rect 12341 13018 12407 13021
rect 8845 13016 12407 13018
rect 8845 12960 8850 13016
rect 8906 12960 12346 13016
rect 12402 12960 12407 13016
rect 8845 12958 12407 12960
rect 8845 12955 8911 12958
rect 12341 12955 12407 12958
rect 9857 12746 9923 12749
rect 17401 12746 17467 12749
rect 9857 12744 17467 12746
rect 9857 12688 9862 12744
rect 9918 12688 17406 12744
rect 17462 12688 17467 12744
rect 9857 12686 17467 12688
rect 9857 12683 9923 12686
rect 17401 12683 17467 12686
rect 9121 12610 9187 12613
rect 9397 12610 9463 12613
rect 9121 12608 9463 12610
rect 9121 12552 9126 12608
rect 9182 12552 9402 12608
rect 9458 12552 9463 12608
rect 9121 12550 9463 12552
rect 9121 12547 9187 12550
rect 9397 12547 9463 12550
rect 14457 12610 14523 12613
rect 15193 12610 15259 12613
rect 14457 12608 15259 12610
rect 14457 12552 14462 12608
rect 14518 12552 15198 12608
rect 15254 12552 15259 12608
rect 14457 12550 15259 12552
rect 14457 12547 14523 12550
rect 15193 12547 15259 12550
rect 4332 12544 4652 12545
rect 4332 12480 4340 12544
rect 4404 12480 4420 12544
rect 4484 12480 4500 12544
rect 4564 12480 4580 12544
rect 4644 12480 4652 12544
rect 4332 12479 4652 12480
rect 11110 12544 11430 12545
rect 11110 12480 11118 12544
rect 11182 12480 11198 12544
rect 11262 12480 11278 12544
rect 11342 12480 11358 12544
rect 11422 12480 11430 12544
rect 11110 12479 11430 12480
rect 17887 12544 18207 12545
rect 17887 12480 17895 12544
rect 17959 12480 17975 12544
rect 18039 12480 18055 12544
rect 18119 12480 18135 12544
rect 18199 12480 18207 12544
rect 17887 12479 18207 12480
rect 8150 12412 8156 12476
rect 8220 12474 8226 12476
rect 9121 12474 9187 12477
rect 8220 12472 9187 12474
rect 8220 12416 9126 12472
rect 9182 12416 9187 12472
rect 8220 12414 9187 12416
rect 8220 12412 8226 12414
rect 9121 12411 9187 12414
rect 12433 12474 12499 12477
rect 14549 12474 14615 12477
rect 12433 12472 14615 12474
rect 12433 12416 12438 12472
rect 12494 12416 14554 12472
rect 14610 12416 14615 12472
rect 12433 12414 14615 12416
rect 12433 12411 12499 12414
rect 14549 12411 14615 12414
rect 0 12338 800 12368
rect 1853 12338 1919 12341
rect 0 12336 1919 12338
rect 0 12280 1858 12336
rect 1914 12280 1919 12336
rect 0 12278 1919 12280
rect 0 12248 800 12278
rect 1853 12275 1919 12278
rect 3969 12338 4035 12341
rect 9489 12338 9555 12341
rect 3969 12336 9555 12338
rect 3969 12280 3974 12336
rect 4030 12280 9494 12336
rect 9550 12280 9555 12336
rect 3969 12278 9555 12280
rect 3969 12275 4035 12278
rect 9489 12275 9555 12278
rect 11697 12338 11763 12341
rect 17677 12338 17743 12341
rect 11697 12336 17743 12338
rect 11697 12280 11702 12336
rect 11758 12280 17682 12336
rect 17738 12280 17743 12336
rect 11697 12278 17743 12280
rect 11697 12275 11763 12278
rect 17677 12275 17743 12278
rect 20713 12338 20779 12341
rect 21767 12338 22567 12368
rect 20713 12336 22567 12338
rect 20713 12280 20718 12336
rect 20774 12280 22567 12336
rect 20713 12278 22567 12280
rect 20713 12275 20779 12278
rect 21767 12248 22567 12278
rect 5993 12202 6059 12205
rect 6545 12202 6611 12205
rect 8293 12202 8359 12205
rect 5993 12200 8359 12202
rect 5993 12144 5998 12200
rect 6054 12144 6550 12200
rect 6606 12144 8298 12200
rect 8354 12144 8359 12200
rect 5993 12142 8359 12144
rect 5993 12139 6059 12142
rect 6545 12139 6611 12142
rect 8293 12139 8359 12142
rect 10317 12202 10383 12205
rect 17401 12202 17467 12205
rect 18413 12202 18479 12205
rect 10317 12200 18479 12202
rect 10317 12144 10322 12200
rect 10378 12144 17406 12200
rect 17462 12144 18418 12200
rect 18474 12144 18479 12200
rect 10317 12142 18479 12144
rect 10317 12139 10383 12142
rect 17401 12139 17467 12142
rect 18413 12139 18479 12142
rect 7721 12000 8041 12001
rect 7721 11936 7729 12000
rect 7793 11936 7809 12000
rect 7873 11936 7889 12000
rect 7953 11936 7969 12000
rect 8033 11936 8041 12000
rect 7721 11935 8041 11936
rect 14498 12000 14818 12001
rect 14498 11936 14506 12000
rect 14570 11936 14586 12000
rect 14650 11936 14666 12000
rect 14730 11936 14746 12000
rect 14810 11936 14818 12000
rect 14498 11935 14818 11936
rect 12249 11794 12315 11797
rect 12525 11794 12591 11797
rect 12249 11792 12591 11794
rect 12249 11736 12254 11792
rect 12310 11736 12530 11792
rect 12586 11736 12591 11792
rect 12249 11734 12591 11736
rect 12249 11731 12315 11734
rect 12525 11731 12591 11734
rect 17585 11658 17651 11661
rect 17542 11656 17651 11658
rect 17542 11600 17590 11656
rect 17646 11600 17651 11656
rect 17542 11595 17651 11600
rect 0 11522 800 11552
rect 1577 11522 1643 11525
rect 0 11520 1643 11522
rect 0 11464 1582 11520
rect 1638 11464 1643 11520
rect 0 11462 1643 11464
rect 0 11432 800 11462
rect 1577 11459 1643 11462
rect 12985 11522 13051 11525
rect 16021 11522 16087 11525
rect 12985 11520 16087 11522
rect 12985 11464 12990 11520
rect 13046 11464 16026 11520
rect 16082 11464 16087 11520
rect 12985 11462 16087 11464
rect 12985 11459 13051 11462
rect 16021 11459 16087 11462
rect 17309 11522 17375 11525
rect 17542 11522 17602 11595
rect 17309 11520 17602 11522
rect 17309 11464 17314 11520
rect 17370 11464 17602 11520
rect 17309 11462 17602 11464
rect 19241 11522 19307 11525
rect 21767 11522 22567 11552
rect 19241 11520 22567 11522
rect 19241 11464 19246 11520
rect 19302 11464 22567 11520
rect 19241 11462 22567 11464
rect 17309 11459 17375 11462
rect 19241 11459 19307 11462
rect 4332 11456 4652 11457
rect 4332 11392 4340 11456
rect 4404 11392 4420 11456
rect 4484 11392 4500 11456
rect 4564 11392 4580 11456
rect 4644 11392 4652 11456
rect 4332 11391 4652 11392
rect 11110 11456 11430 11457
rect 11110 11392 11118 11456
rect 11182 11392 11198 11456
rect 11262 11392 11278 11456
rect 11342 11392 11358 11456
rect 11422 11392 11430 11456
rect 11110 11391 11430 11392
rect 17887 11456 18207 11457
rect 17887 11392 17895 11456
rect 17959 11392 17975 11456
rect 18039 11392 18055 11456
rect 18119 11392 18135 11456
rect 18199 11392 18207 11456
rect 21767 11432 22567 11462
rect 17887 11391 18207 11392
rect 14825 11386 14891 11389
rect 15285 11386 15351 11389
rect 14825 11384 15351 11386
rect 14825 11328 14830 11384
rect 14886 11328 15290 11384
rect 15346 11328 15351 11384
rect 14825 11326 15351 11328
rect 14825 11323 14891 11326
rect 15285 11323 15351 11326
rect 7721 10912 8041 10913
rect 7721 10848 7729 10912
rect 7793 10848 7809 10912
rect 7873 10848 7889 10912
rect 7953 10848 7969 10912
rect 8033 10848 8041 10912
rect 7721 10847 8041 10848
rect 14498 10912 14818 10913
rect 14498 10848 14506 10912
rect 14570 10848 14586 10912
rect 14650 10848 14666 10912
rect 14730 10848 14746 10912
rect 14810 10848 14818 10912
rect 14498 10847 14818 10848
rect 18689 10706 18755 10709
rect 21767 10706 22567 10736
rect 18689 10704 22567 10706
rect 18689 10648 18694 10704
rect 18750 10648 22567 10704
rect 18689 10646 22567 10648
rect 18689 10643 18755 10646
rect 21767 10616 22567 10646
rect 6637 10570 6703 10573
rect 7557 10570 7623 10573
rect 6637 10568 7623 10570
rect 6637 10512 6642 10568
rect 6698 10512 7562 10568
rect 7618 10512 7623 10568
rect 6637 10510 7623 10512
rect 6637 10507 6703 10510
rect 7557 10507 7623 10510
rect 0 10434 800 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 800 10374
rect 1577 10371 1643 10374
rect 13077 10434 13143 10437
rect 16389 10434 16455 10437
rect 17217 10434 17283 10437
rect 13077 10432 17283 10434
rect 13077 10376 13082 10432
rect 13138 10376 16394 10432
rect 16450 10376 17222 10432
rect 17278 10376 17283 10432
rect 13077 10374 17283 10376
rect 13077 10371 13143 10374
rect 16389 10371 16455 10374
rect 17217 10371 17283 10374
rect 4332 10368 4652 10369
rect 4332 10304 4340 10368
rect 4404 10304 4420 10368
rect 4484 10304 4500 10368
rect 4564 10304 4580 10368
rect 4644 10304 4652 10368
rect 4332 10303 4652 10304
rect 11110 10368 11430 10369
rect 11110 10304 11118 10368
rect 11182 10304 11198 10368
rect 11262 10304 11278 10368
rect 11342 10304 11358 10368
rect 11422 10304 11430 10368
rect 11110 10303 11430 10304
rect 17887 10368 18207 10369
rect 17887 10304 17895 10368
rect 17959 10304 17975 10368
rect 18039 10304 18055 10368
rect 18119 10304 18135 10368
rect 18199 10304 18207 10368
rect 17887 10303 18207 10304
rect 8293 10298 8359 10301
rect 9949 10298 10015 10301
rect 10409 10298 10475 10301
rect 8293 10296 10475 10298
rect 8293 10240 8298 10296
rect 8354 10240 9954 10296
rect 10010 10240 10414 10296
rect 10470 10240 10475 10296
rect 8293 10238 10475 10240
rect 8293 10235 8359 10238
rect 9949 10235 10015 10238
rect 10409 10235 10475 10238
rect 1209 10162 1275 10165
rect 16665 10162 16731 10165
rect 1209 10160 16731 10162
rect 1209 10104 1214 10160
rect 1270 10104 16670 10160
rect 16726 10104 16731 10160
rect 1209 10102 16731 10104
rect 1209 10099 1275 10102
rect 16665 10099 16731 10102
rect 7373 10026 7439 10029
rect 9489 10026 9555 10029
rect 7373 10024 9555 10026
rect 7373 9968 7378 10024
rect 7434 9968 9494 10024
rect 9550 9968 9555 10024
rect 7373 9966 9555 9968
rect 7373 9963 7439 9966
rect 9489 9963 9555 9966
rect 7721 9824 8041 9825
rect 7721 9760 7729 9824
rect 7793 9760 7809 9824
rect 7873 9760 7889 9824
rect 7953 9760 7969 9824
rect 8033 9760 8041 9824
rect 7721 9759 8041 9760
rect 14498 9824 14818 9825
rect 14498 9760 14506 9824
rect 14570 9760 14586 9824
rect 14650 9760 14666 9824
rect 14730 9760 14746 9824
rect 14810 9760 14818 9824
rect 14498 9759 14818 9760
rect 8937 9754 9003 9757
rect 9489 9754 9555 9757
rect 8937 9752 9555 9754
rect 8937 9696 8942 9752
rect 8998 9696 9494 9752
rect 9550 9696 9555 9752
rect 8937 9694 9555 9696
rect 8937 9691 9003 9694
rect 9489 9691 9555 9694
rect 0 9618 800 9648
rect 1761 9618 1827 9621
rect 0 9616 1827 9618
rect 0 9560 1766 9616
rect 1822 9560 1827 9616
rect 0 9558 1827 9560
rect 0 9528 800 9558
rect 1761 9555 1827 9558
rect 8109 9618 8175 9621
rect 10501 9618 10567 9621
rect 8109 9616 10567 9618
rect 8109 9560 8114 9616
rect 8170 9560 10506 9616
rect 10562 9560 10567 9616
rect 8109 9558 10567 9560
rect 8109 9555 8175 9558
rect 10501 9555 10567 9558
rect 17033 9618 17099 9621
rect 21767 9618 22567 9648
rect 17033 9616 22567 9618
rect 17033 9560 17038 9616
rect 17094 9560 22567 9616
rect 17033 9558 22567 9560
rect 17033 9555 17099 9558
rect 21767 9528 22567 9558
rect 11973 9482 12039 9485
rect 12801 9482 12867 9485
rect 11973 9480 12867 9482
rect 11973 9424 11978 9480
rect 12034 9424 12806 9480
rect 12862 9424 12867 9480
rect 11973 9422 12867 9424
rect 11973 9419 12039 9422
rect 12801 9419 12867 9422
rect 17493 9482 17559 9485
rect 18321 9482 18387 9485
rect 18597 9482 18663 9485
rect 20294 9482 20300 9484
rect 17493 9480 20300 9482
rect 17493 9424 17498 9480
rect 17554 9424 18326 9480
rect 18382 9424 18602 9480
rect 18658 9424 20300 9480
rect 17493 9422 20300 9424
rect 17493 9419 17559 9422
rect 18321 9419 18387 9422
rect 18597 9419 18663 9422
rect 20294 9420 20300 9422
rect 20364 9420 20370 9484
rect 4332 9280 4652 9281
rect 4332 9216 4340 9280
rect 4404 9216 4420 9280
rect 4484 9216 4500 9280
rect 4564 9216 4580 9280
rect 4644 9216 4652 9280
rect 4332 9215 4652 9216
rect 11110 9280 11430 9281
rect 11110 9216 11118 9280
rect 11182 9216 11198 9280
rect 11262 9216 11278 9280
rect 11342 9216 11358 9280
rect 11422 9216 11430 9280
rect 11110 9215 11430 9216
rect 17887 9280 18207 9281
rect 17887 9216 17895 9280
rect 17959 9216 17975 9280
rect 18039 9216 18055 9280
rect 18119 9216 18135 9280
rect 18199 9216 18207 9280
rect 17887 9215 18207 9216
rect 4153 9074 4219 9077
rect 7189 9074 7255 9077
rect 19926 9074 19932 9076
rect 4153 9072 19932 9074
rect 4153 9016 4158 9072
rect 4214 9016 7194 9072
rect 7250 9016 19932 9072
rect 4153 9014 19932 9016
rect 4153 9011 4219 9014
rect 7189 9011 7255 9014
rect 19926 9012 19932 9014
rect 19996 9012 20002 9076
rect 10961 8938 11027 8941
rect 15653 8938 15719 8941
rect 10961 8936 15719 8938
rect 10961 8880 10966 8936
rect 11022 8880 15658 8936
rect 15714 8880 15719 8936
rect 10961 8878 15719 8880
rect 10961 8875 11027 8878
rect 15653 8875 15719 8878
rect 0 8802 800 8832
rect 1945 8802 2011 8805
rect 0 8800 2011 8802
rect 0 8744 1950 8800
rect 2006 8744 2011 8800
rect 0 8742 2011 8744
rect 0 8712 800 8742
rect 1945 8739 2011 8742
rect 20713 8802 20779 8805
rect 21767 8802 22567 8832
rect 20713 8800 22567 8802
rect 20713 8744 20718 8800
rect 20774 8744 22567 8800
rect 20713 8742 22567 8744
rect 20713 8739 20779 8742
rect 7721 8736 8041 8737
rect 7721 8672 7729 8736
rect 7793 8672 7809 8736
rect 7873 8672 7889 8736
rect 7953 8672 7969 8736
rect 8033 8672 8041 8736
rect 7721 8671 8041 8672
rect 14498 8736 14818 8737
rect 14498 8672 14506 8736
rect 14570 8672 14586 8736
rect 14650 8672 14666 8736
rect 14730 8672 14746 8736
rect 14810 8672 14818 8736
rect 21767 8712 22567 8742
rect 14498 8671 14818 8672
rect 12801 8530 12867 8533
rect 16113 8530 16179 8533
rect 12801 8528 16179 8530
rect 12801 8472 12806 8528
rect 12862 8472 16118 8528
rect 16174 8472 16179 8528
rect 12801 8470 16179 8472
rect 12801 8467 12867 8470
rect 16113 8467 16179 8470
rect 18781 8530 18847 8533
rect 19149 8530 19215 8533
rect 18781 8528 19215 8530
rect 18781 8472 18786 8528
rect 18842 8472 19154 8528
rect 19210 8472 19215 8528
rect 18781 8470 19215 8472
rect 18781 8467 18847 8470
rect 19149 8467 19215 8470
rect 1669 8394 1735 8397
rect 15101 8394 15167 8397
rect 19057 8394 19123 8397
rect 1669 8392 15167 8394
rect 1669 8336 1674 8392
rect 1730 8336 15106 8392
rect 15162 8336 15167 8392
rect 1669 8334 15167 8336
rect 1669 8331 1735 8334
rect 15101 8331 15167 8334
rect 15334 8392 19123 8394
rect 15334 8336 19062 8392
rect 19118 8336 19123 8392
rect 15334 8334 19123 8336
rect 14365 8258 14431 8261
rect 15334 8258 15394 8334
rect 19057 8331 19123 8334
rect 14365 8256 15394 8258
rect 14365 8200 14370 8256
rect 14426 8200 15394 8256
rect 14365 8198 15394 8200
rect 14365 8195 14431 8198
rect 4332 8192 4652 8193
rect 4332 8128 4340 8192
rect 4404 8128 4420 8192
rect 4484 8128 4500 8192
rect 4564 8128 4580 8192
rect 4644 8128 4652 8192
rect 4332 8127 4652 8128
rect 11110 8192 11430 8193
rect 11110 8128 11118 8192
rect 11182 8128 11198 8192
rect 11262 8128 11278 8192
rect 11342 8128 11358 8192
rect 11422 8128 11430 8192
rect 11110 8127 11430 8128
rect 17887 8192 18207 8193
rect 17887 8128 17895 8192
rect 17959 8128 17975 8192
rect 18039 8128 18055 8192
rect 18119 8128 18135 8192
rect 18199 8128 18207 8192
rect 17887 8127 18207 8128
rect 0 7986 800 8016
rect 1669 7986 1735 7989
rect 0 7984 1735 7986
rect 0 7928 1674 7984
rect 1730 7928 1735 7984
rect 0 7926 1735 7928
rect 0 7896 800 7926
rect 1669 7923 1735 7926
rect 3509 7986 3575 7989
rect 7833 7986 7899 7989
rect 3509 7984 7899 7986
rect 3509 7928 3514 7984
rect 3570 7928 7838 7984
rect 7894 7928 7899 7984
rect 3509 7926 7899 7928
rect 3509 7923 3575 7926
rect 7833 7923 7899 7926
rect 11237 7986 11303 7989
rect 14917 7986 14983 7989
rect 11237 7984 14983 7986
rect 11237 7928 11242 7984
rect 11298 7928 14922 7984
rect 14978 7928 14983 7984
rect 11237 7926 14983 7928
rect 11237 7923 11303 7926
rect 14917 7923 14983 7926
rect 17953 7986 18019 7989
rect 21767 7986 22567 8016
rect 17953 7984 22567 7986
rect 17953 7928 17958 7984
rect 18014 7928 22567 7984
rect 17953 7926 22567 7928
rect 17953 7923 18019 7926
rect 21767 7896 22567 7926
rect 3693 7850 3759 7853
rect 11697 7850 11763 7853
rect 3693 7848 11763 7850
rect 3693 7792 3698 7848
rect 3754 7792 11702 7848
rect 11758 7792 11763 7848
rect 3693 7790 11763 7792
rect 3693 7787 3759 7790
rect 11697 7787 11763 7790
rect 7721 7648 8041 7649
rect 7721 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7889 7648
rect 7953 7584 7969 7648
rect 8033 7584 8041 7648
rect 7721 7583 8041 7584
rect 14498 7648 14818 7649
rect 14498 7584 14506 7648
rect 14570 7584 14586 7648
rect 14650 7584 14666 7648
rect 14730 7584 14746 7648
rect 14810 7584 14818 7648
rect 14498 7583 14818 7584
rect 9949 7578 10015 7581
rect 12249 7578 12315 7581
rect 9949 7576 12315 7578
rect 9949 7520 9954 7576
rect 10010 7520 12254 7576
rect 12310 7520 12315 7576
rect 9949 7518 12315 7520
rect 9949 7515 10015 7518
rect 12249 7515 12315 7518
rect 12617 7578 12683 7581
rect 13905 7578 13971 7581
rect 12617 7576 13971 7578
rect 12617 7520 12622 7576
rect 12678 7520 13910 7576
rect 13966 7520 13971 7576
rect 12617 7518 13971 7520
rect 12617 7515 12683 7518
rect 13905 7515 13971 7518
rect 17493 7578 17559 7581
rect 18137 7578 18203 7581
rect 17493 7576 18203 7578
rect 17493 7520 17498 7576
rect 17554 7520 18142 7576
rect 18198 7520 18203 7576
rect 17493 7518 18203 7520
rect 17493 7515 17559 7518
rect 18137 7515 18203 7518
rect 8293 7442 8359 7445
rect 20478 7442 20484 7444
rect 8293 7440 20484 7442
rect 8293 7384 8298 7440
rect 8354 7384 20484 7440
rect 8293 7382 20484 7384
rect 8293 7379 8359 7382
rect 20478 7380 20484 7382
rect 20548 7380 20554 7444
rect 11145 7306 11211 7309
rect 16205 7306 16271 7309
rect 11145 7304 16271 7306
rect 11145 7248 11150 7304
rect 11206 7248 16210 7304
rect 16266 7248 16271 7304
rect 11145 7246 16271 7248
rect 11145 7243 11211 7246
rect 16205 7243 16271 7246
rect 16481 7306 16547 7309
rect 17125 7306 17191 7309
rect 16481 7304 17191 7306
rect 16481 7248 16486 7304
rect 16542 7248 17130 7304
rect 17186 7248 17191 7304
rect 16481 7246 17191 7248
rect 16481 7243 16547 7246
rect 17125 7243 17191 7246
rect 20529 7170 20595 7173
rect 21767 7170 22567 7200
rect 20529 7168 22567 7170
rect 20529 7112 20534 7168
rect 20590 7112 22567 7168
rect 20529 7110 22567 7112
rect 20529 7107 20595 7110
rect 4332 7104 4652 7105
rect 4332 7040 4340 7104
rect 4404 7040 4420 7104
rect 4484 7040 4500 7104
rect 4564 7040 4580 7104
rect 4644 7040 4652 7104
rect 4332 7039 4652 7040
rect 11110 7104 11430 7105
rect 11110 7040 11118 7104
rect 11182 7040 11198 7104
rect 11262 7040 11278 7104
rect 11342 7040 11358 7104
rect 11422 7040 11430 7104
rect 11110 7039 11430 7040
rect 17887 7104 18207 7105
rect 17887 7040 17895 7104
rect 17959 7040 17975 7104
rect 18039 7040 18055 7104
rect 18119 7040 18135 7104
rect 18199 7040 18207 7104
rect 21767 7080 22567 7110
rect 17887 7039 18207 7040
rect 7281 7034 7347 7037
rect 8150 7034 8156 7036
rect 7281 7032 8156 7034
rect 7281 6976 7286 7032
rect 7342 6976 8156 7032
rect 7281 6974 8156 6976
rect 7281 6971 7347 6974
rect 8150 6972 8156 6974
rect 8220 6972 8226 7036
rect 0 6898 800 6928
rect 1853 6898 1919 6901
rect 0 6896 1919 6898
rect 0 6840 1858 6896
rect 1914 6840 1919 6896
rect 0 6838 1919 6840
rect 0 6808 800 6838
rect 1853 6835 1919 6838
rect 2221 6898 2287 6901
rect 9121 6898 9187 6901
rect 16573 6898 16639 6901
rect 2221 6896 2790 6898
rect 2221 6840 2226 6896
rect 2282 6840 2790 6896
rect 2221 6838 2790 6840
rect 2221 6835 2287 6838
rect 2730 6762 2790 6838
rect 9121 6896 16639 6898
rect 9121 6840 9126 6896
rect 9182 6840 16578 6896
rect 16634 6840 16639 6896
rect 9121 6838 16639 6840
rect 9121 6835 9187 6838
rect 16573 6835 16639 6838
rect 15377 6762 15443 6765
rect 15745 6762 15811 6765
rect 2730 6760 15811 6762
rect 2730 6704 15382 6760
rect 15438 6704 15750 6760
rect 15806 6704 15811 6760
rect 2730 6702 15811 6704
rect 15377 6699 15443 6702
rect 15745 6699 15811 6702
rect 17033 6762 17099 6765
rect 18321 6762 18387 6765
rect 18781 6762 18847 6765
rect 17033 6760 18847 6762
rect 17033 6704 17038 6760
rect 17094 6704 18326 6760
rect 18382 6704 18786 6760
rect 18842 6704 18847 6760
rect 17033 6702 18847 6704
rect 17033 6699 17099 6702
rect 18321 6699 18387 6702
rect 18781 6699 18847 6702
rect 1761 6626 1827 6629
rect 5349 6626 5415 6629
rect 1761 6624 5415 6626
rect 1761 6568 1766 6624
rect 1822 6568 5354 6624
rect 5410 6568 5415 6624
rect 1761 6566 5415 6568
rect 1761 6563 1827 6566
rect 5349 6563 5415 6566
rect 11605 6626 11671 6629
rect 12341 6626 12407 6629
rect 11605 6624 12407 6626
rect 11605 6568 11610 6624
rect 11666 6568 12346 6624
rect 12402 6568 12407 6624
rect 11605 6566 12407 6568
rect 11605 6563 11671 6566
rect 12341 6563 12407 6566
rect 15653 6626 15719 6629
rect 17309 6626 17375 6629
rect 15653 6624 17375 6626
rect 15653 6568 15658 6624
rect 15714 6568 17314 6624
rect 17370 6568 17375 6624
rect 15653 6566 17375 6568
rect 15653 6563 15719 6566
rect 17309 6563 17375 6566
rect 7721 6560 8041 6561
rect 7721 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7889 6560
rect 7953 6496 7969 6560
rect 8033 6496 8041 6560
rect 7721 6495 8041 6496
rect 14498 6560 14818 6561
rect 14498 6496 14506 6560
rect 14570 6496 14586 6560
rect 14650 6496 14666 6560
rect 14730 6496 14746 6560
rect 14810 6496 14818 6560
rect 14498 6495 14818 6496
rect 7465 6354 7531 6357
rect 7054 6352 7531 6354
rect 7054 6296 7470 6352
rect 7526 6296 7531 6352
rect 7054 6294 7531 6296
rect 7054 6221 7114 6294
rect 7465 6291 7531 6294
rect 7005 6216 7114 6221
rect 7005 6160 7010 6216
rect 7066 6160 7114 6216
rect 7005 6158 7114 6160
rect 7465 6218 7531 6221
rect 18873 6218 18939 6221
rect 7465 6216 18939 6218
rect 7465 6160 7470 6216
rect 7526 6160 18878 6216
rect 18934 6160 18939 6216
rect 7465 6158 18939 6160
rect 7005 6155 7071 6158
rect 7465 6155 7531 6158
rect 18873 6155 18939 6158
rect 0 6082 800 6112
rect 1945 6082 2011 6085
rect 0 6080 2011 6082
rect 0 6024 1950 6080
rect 2006 6024 2011 6080
rect 0 6022 2011 6024
rect 0 5992 800 6022
rect 1945 6019 2011 6022
rect 19241 6082 19307 6085
rect 21767 6082 22567 6112
rect 19241 6080 22567 6082
rect 19241 6024 19246 6080
rect 19302 6024 22567 6080
rect 19241 6022 22567 6024
rect 19241 6019 19307 6022
rect 4332 6016 4652 6017
rect 4332 5952 4340 6016
rect 4404 5952 4420 6016
rect 4484 5952 4500 6016
rect 4564 5952 4580 6016
rect 4644 5952 4652 6016
rect 4332 5951 4652 5952
rect 11110 6016 11430 6017
rect 11110 5952 11118 6016
rect 11182 5952 11198 6016
rect 11262 5952 11278 6016
rect 11342 5952 11358 6016
rect 11422 5952 11430 6016
rect 11110 5951 11430 5952
rect 17887 6016 18207 6017
rect 17887 5952 17895 6016
rect 17959 5952 17975 6016
rect 18039 5952 18055 6016
rect 18119 5952 18135 6016
rect 18199 5952 18207 6016
rect 21767 5992 22567 6022
rect 17887 5951 18207 5952
rect 19977 5946 20043 5949
rect 20110 5946 20116 5948
rect 19977 5944 20116 5946
rect 19977 5888 19982 5944
rect 20038 5888 20116 5944
rect 19977 5886 20116 5888
rect 19977 5883 20043 5886
rect 20110 5884 20116 5886
rect 20180 5884 20186 5948
rect 6361 5810 6427 5813
rect 19333 5810 19399 5813
rect 6361 5808 19399 5810
rect 6361 5752 6366 5808
rect 6422 5752 19338 5808
rect 19394 5752 19399 5808
rect 6361 5750 19399 5752
rect 6361 5747 6427 5750
rect 19333 5747 19399 5750
rect 1853 5674 1919 5677
rect 17677 5674 17743 5677
rect 1853 5672 17743 5674
rect 1853 5616 1858 5672
rect 1914 5616 17682 5672
rect 17738 5616 17743 5672
rect 1853 5614 17743 5616
rect 1853 5611 1919 5614
rect 17677 5611 17743 5614
rect 9029 5538 9095 5541
rect 9489 5538 9555 5541
rect 9029 5536 9555 5538
rect 9029 5480 9034 5536
rect 9090 5480 9494 5536
rect 9550 5480 9555 5536
rect 9029 5478 9555 5480
rect 9029 5475 9095 5478
rect 9489 5475 9555 5478
rect 7721 5472 8041 5473
rect 7721 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7889 5472
rect 7953 5408 7969 5472
rect 8033 5408 8041 5472
rect 7721 5407 8041 5408
rect 14498 5472 14818 5473
rect 14498 5408 14506 5472
rect 14570 5408 14586 5472
rect 14650 5408 14666 5472
rect 14730 5408 14746 5472
rect 14810 5408 14818 5472
rect 14498 5407 14818 5408
rect 9438 5340 9444 5404
rect 9508 5402 9514 5404
rect 9581 5402 9647 5405
rect 9508 5400 9647 5402
rect 9508 5344 9586 5400
rect 9642 5344 9647 5400
rect 9508 5342 9647 5344
rect 9508 5340 9514 5342
rect 9581 5339 9647 5342
rect 0 5266 800 5296
rect 2037 5266 2103 5269
rect 0 5264 2103 5266
rect 0 5208 2042 5264
rect 2098 5208 2103 5264
rect 0 5206 2103 5208
rect 0 5176 800 5206
rect 2037 5203 2103 5206
rect 9305 5266 9371 5269
rect 14733 5266 14799 5269
rect 9305 5264 9506 5266
rect 9305 5208 9310 5264
rect 9366 5208 9506 5264
rect 9305 5206 9506 5208
rect 9305 5203 9371 5206
rect 9446 5130 9506 5206
rect 13678 5264 14799 5266
rect 13678 5208 14738 5264
rect 14794 5208 14799 5264
rect 13678 5206 14799 5208
rect 9581 5130 9647 5133
rect 9446 5128 9647 5130
rect 9446 5072 9586 5128
rect 9642 5072 9647 5128
rect 9446 5070 9647 5072
rect 9581 5067 9647 5070
rect 9857 5130 9923 5133
rect 12893 5130 12959 5133
rect 13678 5130 13738 5206
rect 14733 5203 14799 5206
rect 20529 5266 20595 5269
rect 21767 5266 22567 5296
rect 20529 5264 22567 5266
rect 20529 5208 20534 5264
rect 20590 5208 22567 5264
rect 20529 5206 22567 5208
rect 20529 5203 20595 5206
rect 21767 5176 22567 5206
rect 9857 5128 13738 5130
rect 9857 5072 9862 5128
rect 9918 5072 12898 5128
rect 12954 5072 13738 5128
rect 9857 5070 13738 5072
rect 13813 5130 13879 5133
rect 17493 5130 17559 5133
rect 13813 5128 17559 5130
rect 13813 5072 13818 5128
rect 13874 5072 17498 5128
rect 17554 5072 17559 5128
rect 13813 5070 17559 5072
rect 9857 5067 9923 5070
rect 12893 5067 12959 5070
rect 13813 5067 13879 5070
rect 17493 5067 17559 5070
rect 4332 4928 4652 4929
rect 4332 4864 4340 4928
rect 4404 4864 4420 4928
rect 4484 4864 4500 4928
rect 4564 4864 4580 4928
rect 4644 4864 4652 4928
rect 4332 4863 4652 4864
rect 11110 4928 11430 4929
rect 11110 4864 11118 4928
rect 11182 4864 11198 4928
rect 11262 4864 11278 4928
rect 11342 4864 11358 4928
rect 11422 4864 11430 4928
rect 11110 4863 11430 4864
rect 17887 4928 18207 4929
rect 17887 4864 17895 4928
rect 17959 4864 17975 4928
rect 18039 4864 18055 4928
rect 18119 4864 18135 4928
rect 18199 4864 18207 4928
rect 17887 4863 18207 4864
rect 9213 4858 9279 4861
rect 9438 4858 9444 4860
rect 9213 4856 9444 4858
rect 9213 4800 9218 4856
rect 9274 4800 9444 4856
rect 9213 4798 9444 4800
rect 9213 4795 9279 4798
rect 9438 4796 9444 4798
rect 9508 4858 9514 4860
rect 9581 4858 9647 4861
rect 9508 4856 9647 4858
rect 9508 4800 9586 4856
rect 9642 4800 9647 4856
rect 9508 4798 9647 4800
rect 9508 4796 9514 4798
rect 9581 4795 9647 4798
rect 7097 4586 7163 4589
rect 7097 4584 12450 4586
rect 7097 4528 7102 4584
rect 7158 4528 12450 4584
rect 7097 4526 12450 4528
rect 7097 4523 7163 4526
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 7721 4384 8041 4385
rect 7721 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7889 4384
rect 7953 4320 7969 4384
rect 8033 4320 8041 4384
rect 7721 4319 8041 4320
rect 12390 4178 12450 4526
rect 20713 4450 20779 4453
rect 21767 4450 22567 4480
rect 20713 4448 22567 4450
rect 20713 4392 20718 4448
rect 20774 4392 22567 4448
rect 20713 4390 22567 4392
rect 20713 4387 20779 4390
rect 14498 4384 14818 4385
rect 14498 4320 14506 4384
rect 14570 4320 14586 4384
rect 14650 4320 14666 4384
rect 14730 4320 14746 4384
rect 14810 4320 14818 4384
rect 21767 4360 22567 4390
rect 14498 4319 14818 4320
rect 20253 4178 20319 4181
rect 12390 4176 20319 4178
rect 12390 4120 20258 4176
rect 20314 4120 20319 4176
rect 12390 4118 20319 4120
rect 20253 4115 20319 4118
rect 4332 3840 4652 3841
rect 4332 3776 4340 3840
rect 4404 3776 4420 3840
rect 4484 3776 4500 3840
rect 4564 3776 4580 3840
rect 4644 3776 4652 3840
rect 4332 3775 4652 3776
rect 11110 3840 11430 3841
rect 11110 3776 11118 3840
rect 11182 3776 11198 3840
rect 11262 3776 11278 3840
rect 11342 3776 11358 3840
rect 11422 3776 11430 3840
rect 11110 3775 11430 3776
rect 17887 3840 18207 3841
rect 17887 3776 17895 3840
rect 17959 3776 17975 3840
rect 18039 3776 18055 3840
rect 18119 3776 18135 3840
rect 18199 3776 18207 3840
rect 17887 3775 18207 3776
rect 3233 3634 3299 3637
rect 4521 3634 4587 3637
rect 3233 3632 4587 3634
rect 3233 3576 3238 3632
rect 3294 3576 4526 3632
rect 4582 3576 4587 3632
rect 3233 3574 4587 3576
rect 3233 3571 3299 3574
rect 4521 3571 4587 3574
rect 9673 3634 9739 3637
rect 13905 3634 13971 3637
rect 9673 3632 13971 3634
rect 9673 3576 9678 3632
rect 9734 3576 13910 3632
rect 13966 3576 13971 3632
rect 9673 3574 13971 3576
rect 9673 3571 9739 3574
rect 13905 3571 13971 3574
rect 17953 3634 18019 3637
rect 21767 3634 22567 3664
rect 17953 3632 22567 3634
rect 17953 3576 17958 3632
rect 18014 3576 22567 3632
rect 17953 3574 22567 3576
rect 17953 3571 18019 3574
rect 21767 3544 22567 3574
rect 8150 3436 8156 3500
rect 8220 3498 8226 3500
rect 19517 3498 19583 3501
rect 8220 3496 19583 3498
rect 8220 3440 19522 3496
rect 19578 3440 19583 3496
rect 8220 3438 19583 3440
rect 8220 3436 8226 3438
rect 19517 3435 19583 3438
rect 0 3362 800 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 800 3302
rect 3969 3299 4035 3302
rect 15377 3362 15443 3365
rect 18137 3362 18203 3365
rect 15377 3360 18203 3362
rect 15377 3304 15382 3360
rect 15438 3304 18142 3360
rect 18198 3304 18203 3360
rect 15377 3302 18203 3304
rect 15377 3299 15443 3302
rect 18137 3299 18203 3302
rect 7721 3296 8041 3297
rect 7721 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7889 3296
rect 7953 3232 7969 3296
rect 8033 3232 8041 3296
rect 7721 3231 8041 3232
rect 14498 3296 14818 3297
rect 14498 3232 14506 3296
rect 14570 3232 14586 3296
rect 14650 3232 14666 3296
rect 14730 3232 14746 3296
rect 14810 3232 14818 3296
rect 14498 3231 14818 3232
rect 12433 3226 12499 3229
rect 12893 3226 12959 3229
rect 12433 3224 12959 3226
rect 12433 3168 12438 3224
rect 12494 3168 12898 3224
rect 12954 3168 12959 3224
rect 12433 3166 12959 3168
rect 12433 3163 12499 3166
rect 12893 3163 12959 3166
rect 4332 2752 4652 2753
rect 4332 2688 4340 2752
rect 4404 2688 4420 2752
rect 4484 2688 4500 2752
rect 4564 2688 4580 2752
rect 4644 2688 4652 2752
rect 4332 2687 4652 2688
rect 11110 2752 11430 2753
rect 11110 2688 11118 2752
rect 11182 2688 11198 2752
rect 11262 2688 11278 2752
rect 11342 2688 11358 2752
rect 11422 2688 11430 2752
rect 11110 2687 11430 2688
rect 17887 2752 18207 2753
rect 17887 2688 17895 2752
rect 17959 2688 17975 2752
rect 18039 2688 18055 2752
rect 18119 2688 18135 2752
rect 18199 2688 18207 2752
rect 17887 2687 18207 2688
rect 0 2546 800 2576
rect 2773 2546 2839 2549
rect 0 2544 2839 2546
rect 0 2488 2778 2544
rect 2834 2488 2839 2544
rect 0 2486 2839 2488
rect 0 2456 800 2486
rect 2773 2483 2839 2486
rect 18873 2546 18939 2549
rect 21767 2546 22567 2576
rect 18873 2544 22567 2546
rect 18873 2488 18878 2544
rect 18934 2488 22567 2544
rect 18873 2486 22567 2488
rect 18873 2483 18939 2486
rect 21767 2456 22567 2486
rect 7721 2208 8041 2209
rect 7721 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7889 2208
rect 7953 2144 7969 2208
rect 8033 2144 8041 2208
rect 7721 2143 8041 2144
rect 14498 2208 14818 2209
rect 14498 2144 14506 2208
rect 14570 2144 14586 2208
rect 14650 2144 14666 2208
rect 14730 2144 14746 2208
rect 14810 2144 14818 2208
rect 14498 2143 14818 2144
rect 0 1730 800 1760
rect 2865 1730 2931 1733
rect 0 1728 2931 1730
rect 0 1672 2870 1728
rect 2926 1672 2931 1728
rect 0 1670 2931 1672
rect 0 1640 800 1670
rect 2865 1667 2931 1670
rect 19977 1730 20043 1733
rect 21767 1730 22567 1760
rect 19977 1728 22567 1730
rect 19977 1672 19982 1728
rect 20038 1672 22567 1728
rect 19977 1670 22567 1672
rect 19977 1667 20043 1670
rect 21767 1640 22567 1670
rect 0 914 800 944
rect 1853 914 1919 917
rect 0 912 1919 914
rect 0 856 1858 912
rect 1914 856 1919 912
rect 0 854 1919 856
rect 0 824 800 854
rect 1853 851 1919 854
rect 17585 914 17651 917
rect 21767 914 22567 944
rect 17585 912 22567 914
rect 17585 856 17590 912
rect 17646 856 22567 912
rect 17585 854 22567 856
rect 17585 851 17651 854
rect 21767 824 22567 854
rect 16941 98 17007 101
rect 21767 98 22567 128
rect 16941 96 22567 98
rect 16941 40 16946 96
rect 17002 40 22567 96
rect 16941 38 22567 40
rect 16941 35 17007 38
rect 21767 8 22567 38
<< via3 >>
rect 4340 22332 4404 22336
rect 4340 22276 4344 22332
rect 4344 22276 4400 22332
rect 4400 22276 4404 22332
rect 4340 22272 4404 22276
rect 4420 22332 4484 22336
rect 4420 22276 4424 22332
rect 4424 22276 4480 22332
rect 4480 22276 4484 22332
rect 4420 22272 4484 22276
rect 4500 22332 4564 22336
rect 4500 22276 4504 22332
rect 4504 22276 4560 22332
rect 4560 22276 4564 22332
rect 4500 22272 4564 22276
rect 4580 22332 4644 22336
rect 4580 22276 4584 22332
rect 4584 22276 4640 22332
rect 4640 22276 4644 22332
rect 4580 22272 4644 22276
rect 11118 22332 11182 22336
rect 11118 22276 11122 22332
rect 11122 22276 11178 22332
rect 11178 22276 11182 22332
rect 11118 22272 11182 22276
rect 11198 22332 11262 22336
rect 11198 22276 11202 22332
rect 11202 22276 11258 22332
rect 11258 22276 11262 22332
rect 11198 22272 11262 22276
rect 11278 22332 11342 22336
rect 11278 22276 11282 22332
rect 11282 22276 11338 22332
rect 11338 22276 11342 22332
rect 11278 22272 11342 22276
rect 11358 22332 11422 22336
rect 11358 22276 11362 22332
rect 11362 22276 11418 22332
rect 11418 22276 11422 22332
rect 11358 22272 11422 22276
rect 17895 22332 17959 22336
rect 17895 22276 17899 22332
rect 17899 22276 17955 22332
rect 17955 22276 17959 22332
rect 17895 22272 17959 22276
rect 17975 22332 18039 22336
rect 17975 22276 17979 22332
rect 17979 22276 18035 22332
rect 18035 22276 18039 22332
rect 17975 22272 18039 22276
rect 18055 22332 18119 22336
rect 18055 22276 18059 22332
rect 18059 22276 18115 22332
rect 18115 22276 18119 22332
rect 18055 22272 18119 22276
rect 18135 22332 18199 22336
rect 18135 22276 18139 22332
rect 18139 22276 18195 22332
rect 18195 22276 18199 22332
rect 18135 22272 18199 22276
rect 7729 21788 7793 21792
rect 7729 21732 7733 21788
rect 7733 21732 7789 21788
rect 7789 21732 7793 21788
rect 7729 21728 7793 21732
rect 7809 21788 7873 21792
rect 7809 21732 7813 21788
rect 7813 21732 7869 21788
rect 7869 21732 7873 21788
rect 7809 21728 7873 21732
rect 7889 21788 7953 21792
rect 7889 21732 7893 21788
rect 7893 21732 7949 21788
rect 7949 21732 7953 21788
rect 7889 21728 7953 21732
rect 7969 21788 8033 21792
rect 7969 21732 7973 21788
rect 7973 21732 8029 21788
rect 8029 21732 8033 21788
rect 7969 21728 8033 21732
rect 14506 21788 14570 21792
rect 14506 21732 14510 21788
rect 14510 21732 14566 21788
rect 14566 21732 14570 21788
rect 14506 21728 14570 21732
rect 14586 21788 14650 21792
rect 14586 21732 14590 21788
rect 14590 21732 14646 21788
rect 14646 21732 14650 21788
rect 14586 21728 14650 21732
rect 14666 21788 14730 21792
rect 14666 21732 14670 21788
rect 14670 21732 14726 21788
rect 14726 21732 14730 21788
rect 14666 21728 14730 21732
rect 14746 21788 14810 21792
rect 14746 21732 14750 21788
rect 14750 21732 14806 21788
rect 14806 21732 14810 21788
rect 14746 21728 14810 21732
rect 4340 21244 4404 21248
rect 4340 21188 4344 21244
rect 4344 21188 4400 21244
rect 4400 21188 4404 21244
rect 4340 21184 4404 21188
rect 4420 21244 4484 21248
rect 4420 21188 4424 21244
rect 4424 21188 4480 21244
rect 4480 21188 4484 21244
rect 4420 21184 4484 21188
rect 4500 21244 4564 21248
rect 4500 21188 4504 21244
rect 4504 21188 4560 21244
rect 4560 21188 4564 21244
rect 4500 21184 4564 21188
rect 4580 21244 4644 21248
rect 4580 21188 4584 21244
rect 4584 21188 4640 21244
rect 4640 21188 4644 21244
rect 4580 21184 4644 21188
rect 11118 21244 11182 21248
rect 11118 21188 11122 21244
rect 11122 21188 11178 21244
rect 11178 21188 11182 21244
rect 11118 21184 11182 21188
rect 11198 21244 11262 21248
rect 11198 21188 11202 21244
rect 11202 21188 11258 21244
rect 11258 21188 11262 21244
rect 11198 21184 11262 21188
rect 11278 21244 11342 21248
rect 11278 21188 11282 21244
rect 11282 21188 11338 21244
rect 11338 21188 11342 21244
rect 11278 21184 11342 21188
rect 11358 21244 11422 21248
rect 11358 21188 11362 21244
rect 11362 21188 11418 21244
rect 11418 21188 11422 21244
rect 11358 21184 11422 21188
rect 17895 21244 17959 21248
rect 17895 21188 17899 21244
rect 17899 21188 17955 21244
rect 17955 21188 17959 21244
rect 17895 21184 17959 21188
rect 17975 21244 18039 21248
rect 17975 21188 17979 21244
rect 17979 21188 18035 21244
rect 18035 21188 18039 21244
rect 17975 21184 18039 21188
rect 18055 21244 18119 21248
rect 18055 21188 18059 21244
rect 18059 21188 18115 21244
rect 18115 21188 18119 21244
rect 18055 21184 18119 21188
rect 18135 21244 18199 21248
rect 18135 21188 18139 21244
rect 18139 21188 18195 21244
rect 18195 21188 18199 21244
rect 18135 21184 18199 21188
rect 20300 20708 20364 20772
rect 20484 20708 20548 20772
rect 7729 20700 7793 20704
rect 7729 20644 7733 20700
rect 7733 20644 7789 20700
rect 7789 20644 7793 20700
rect 7729 20640 7793 20644
rect 7809 20700 7873 20704
rect 7809 20644 7813 20700
rect 7813 20644 7869 20700
rect 7869 20644 7873 20700
rect 7809 20640 7873 20644
rect 7889 20700 7953 20704
rect 7889 20644 7893 20700
rect 7893 20644 7949 20700
rect 7949 20644 7953 20700
rect 7889 20640 7953 20644
rect 7969 20700 8033 20704
rect 7969 20644 7973 20700
rect 7973 20644 8029 20700
rect 8029 20644 8033 20700
rect 7969 20640 8033 20644
rect 14506 20700 14570 20704
rect 14506 20644 14510 20700
rect 14510 20644 14566 20700
rect 14566 20644 14570 20700
rect 14506 20640 14570 20644
rect 14586 20700 14650 20704
rect 14586 20644 14590 20700
rect 14590 20644 14646 20700
rect 14646 20644 14650 20700
rect 14586 20640 14650 20644
rect 14666 20700 14730 20704
rect 14666 20644 14670 20700
rect 14670 20644 14726 20700
rect 14726 20644 14730 20700
rect 14666 20640 14730 20644
rect 14746 20700 14810 20704
rect 14746 20644 14750 20700
rect 14750 20644 14806 20700
rect 14806 20644 14810 20700
rect 14746 20640 14810 20644
rect 4340 20156 4404 20160
rect 4340 20100 4344 20156
rect 4344 20100 4400 20156
rect 4400 20100 4404 20156
rect 4340 20096 4404 20100
rect 4420 20156 4484 20160
rect 4420 20100 4424 20156
rect 4424 20100 4480 20156
rect 4480 20100 4484 20156
rect 4420 20096 4484 20100
rect 4500 20156 4564 20160
rect 4500 20100 4504 20156
rect 4504 20100 4560 20156
rect 4560 20100 4564 20156
rect 4500 20096 4564 20100
rect 4580 20156 4644 20160
rect 4580 20100 4584 20156
rect 4584 20100 4640 20156
rect 4640 20100 4644 20156
rect 4580 20096 4644 20100
rect 11118 20156 11182 20160
rect 11118 20100 11122 20156
rect 11122 20100 11178 20156
rect 11178 20100 11182 20156
rect 11118 20096 11182 20100
rect 11198 20156 11262 20160
rect 11198 20100 11202 20156
rect 11202 20100 11258 20156
rect 11258 20100 11262 20156
rect 11198 20096 11262 20100
rect 11278 20156 11342 20160
rect 11278 20100 11282 20156
rect 11282 20100 11338 20156
rect 11338 20100 11342 20156
rect 11278 20096 11342 20100
rect 11358 20156 11422 20160
rect 11358 20100 11362 20156
rect 11362 20100 11418 20156
rect 11418 20100 11422 20156
rect 11358 20096 11422 20100
rect 17895 20156 17959 20160
rect 17895 20100 17899 20156
rect 17899 20100 17955 20156
rect 17955 20100 17959 20156
rect 17895 20096 17959 20100
rect 17975 20156 18039 20160
rect 17975 20100 17979 20156
rect 17979 20100 18035 20156
rect 18035 20100 18039 20156
rect 17975 20096 18039 20100
rect 18055 20156 18119 20160
rect 18055 20100 18059 20156
rect 18059 20100 18115 20156
rect 18115 20100 18119 20156
rect 18055 20096 18119 20100
rect 18135 20156 18199 20160
rect 18135 20100 18139 20156
rect 18139 20100 18195 20156
rect 18195 20100 18199 20156
rect 18135 20096 18199 20100
rect 19932 19620 19996 19684
rect 7729 19612 7793 19616
rect 7729 19556 7733 19612
rect 7733 19556 7789 19612
rect 7789 19556 7793 19612
rect 7729 19552 7793 19556
rect 7809 19612 7873 19616
rect 7809 19556 7813 19612
rect 7813 19556 7869 19612
rect 7869 19556 7873 19612
rect 7809 19552 7873 19556
rect 7889 19612 7953 19616
rect 7889 19556 7893 19612
rect 7893 19556 7949 19612
rect 7949 19556 7953 19612
rect 7889 19552 7953 19556
rect 7969 19612 8033 19616
rect 7969 19556 7973 19612
rect 7973 19556 8029 19612
rect 8029 19556 8033 19612
rect 7969 19552 8033 19556
rect 14506 19612 14570 19616
rect 14506 19556 14510 19612
rect 14510 19556 14566 19612
rect 14566 19556 14570 19612
rect 14506 19552 14570 19556
rect 14586 19612 14650 19616
rect 14586 19556 14590 19612
rect 14590 19556 14646 19612
rect 14646 19556 14650 19612
rect 14586 19552 14650 19556
rect 14666 19612 14730 19616
rect 14666 19556 14670 19612
rect 14670 19556 14726 19612
rect 14726 19556 14730 19612
rect 14666 19552 14730 19556
rect 14746 19612 14810 19616
rect 14746 19556 14750 19612
rect 14750 19556 14806 19612
rect 14806 19556 14810 19612
rect 14746 19552 14810 19556
rect 20116 19484 20180 19548
rect 14964 19272 15028 19276
rect 14964 19216 14978 19272
rect 14978 19216 15028 19272
rect 14964 19212 15028 19216
rect 4340 19068 4404 19072
rect 4340 19012 4344 19068
rect 4344 19012 4400 19068
rect 4400 19012 4404 19068
rect 4340 19008 4404 19012
rect 4420 19068 4484 19072
rect 4420 19012 4424 19068
rect 4424 19012 4480 19068
rect 4480 19012 4484 19068
rect 4420 19008 4484 19012
rect 4500 19068 4564 19072
rect 4500 19012 4504 19068
rect 4504 19012 4560 19068
rect 4560 19012 4564 19068
rect 4500 19008 4564 19012
rect 4580 19068 4644 19072
rect 4580 19012 4584 19068
rect 4584 19012 4640 19068
rect 4640 19012 4644 19068
rect 4580 19008 4644 19012
rect 11118 19068 11182 19072
rect 11118 19012 11122 19068
rect 11122 19012 11178 19068
rect 11178 19012 11182 19068
rect 11118 19008 11182 19012
rect 11198 19068 11262 19072
rect 11198 19012 11202 19068
rect 11202 19012 11258 19068
rect 11258 19012 11262 19068
rect 11198 19008 11262 19012
rect 11278 19068 11342 19072
rect 11278 19012 11282 19068
rect 11282 19012 11338 19068
rect 11338 19012 11342 19068
rect 11278 19008 11342 19012
rect 11358 19068 11422 19072
rect 11358 19012 11362 19068
rect 11362 19012 11418 19068
rect 11418 19012 11422 19068
rect 11358 19008 11422 19012
rect 17895 19068 17959 19072
rect 17895 19012 17899 19068
rect 17899 19012 17955 19068
rect 17955 19012 17959 19068
rect 17895 19008 17959 19012
rect 17975 19068 18039 19072
rect 17975 19012 17979 19068
rect 17979 19012 18035 19068
rect 18035 19012 18039 19068
rect 17975 19008 18039 19012
rect 18055 19068 18119 19072
rect 18055 19012 18059 19068
rect 18059 19012 18115 19068
rect 18115 19012 18119 19068
rect 18055 19008 18119 19012
rect 18135 19068 18199 19072
rect 18135 19012 18139 19068
rect 18139 19012 18195 19068
rect 18195 19012 18199 19068
rect 18135 19008 18199 19012
rect 7729 18524 7793 18528
rect 7729 18468 7733 18524
rect 7733 18468 7789 18524
rect 7789 18468 7793 18524
rect 7729 18464 7793 18468
rect 7809 18524 7873 18528
rect 7809 18468 7813 18524
rect 7813 18468 7869 18524
rect 7869 18468 7873 18524
rect 7809 18464 7873 18468
rect 7889 18524 7953 18528
rect 7889 18468 7893 18524
rect 7893 18468 7949 18524
rect 7949 18468 7953 18524
rect 7889 18464 7953 18468
rect 7969 18524 8033 18528
rect 7969 18468 7973 18524
rect 7973 18468 8029 18524
rect 8029 18468 8033 18524
rect 7969 18464 8033 18468
rect 14506 18524 14570 18528
rect 14506 18468 14510 18524
rect 14510 18468 14566 18524
rect 14566 18468 14570 18524
rect 14506 18464 14570 18468
rect 14586 18524 14650 18528
rect 14586 18468 14590 18524
rect 14590 18468 14646 18524
rect 14646 18468 14650 18524
rect 14586 18464 14650 18468
rect 14666 18524 14730 18528
rect 14666 18468 14670 18524
rect 14670 18468 14726 18524
rect 14726 18468 14730 18524
rect 14666 18464 14730 18468
rect 14746 18524 14810 18528
rect 14746 18468 14750 18524
rect 14750 18468 14806 18524
rect 14806 18468 14810 18524
rect 14746 18464 14810 18468
rect 4340 17980 4404 17984
rect 4340 17924 4344 17980
rect 4344 17924 4400 17980
rect 4400 17924 4404 17980
rect 4340 17920 4404 17924
rect 4420 17980 4484 17984
rect 4420 17924 4424 17980
rect 4424 17924 4480 17980
rect 4480 17924 4484 17980
rect 4420 17920 4484 17924
rect 4500 17980 4564 17984
rect 4500 17924 4504 17980
rect 4504 17924 4560 17980
rect 4560 17924 4564 17980
rect 4500 17920 4564 17924
rect 4580 17980 4644 17984
rect 4580 17924 4584 17980
rect 4584 17924 4640 17980
rect 4640 17924 4644 17980
rect 4580 17920 4644 17924
rect 11118 17980 11182 17984
rect 11118 17924 11122 17980
rect 11122 17924 11178 17980
rect 11178 17924 11182 17980
rect 11118 17920 11182 17924
rect 11198 17980 11262 17984
rect 11198 17924 11202 17980
rect 11202 17924 11258 17980
rect 11258 17924 11262 17980
rect 11198 17920 11262 17924
rect 11278 17980 11342 17984
rect 11278 17924 11282 17980
rect 11282 17924 11338 17980
rect 11338 17924 11342 17980
rect 11278 17920 11342 17924
rect 11358 17980 11422 17984
rect 11358 17924 11362 17980
rect 11362 17924 11418 17980
rect 11418 17924 11422 17980
rect 11358 17920 11422 17924
rect 17895 17980 17959 17984
rect 17895 17924 17899 17980
rect 17899 17924 17955 17980
rect 17955 17924 17959 17980
rect 17895 17920 17959 17924
rect 17975 17980 18039 17984
rect 17975 17924 17979 17980
rect 17979 17924 18035 17980
rect 18035 17924 18039 17980
rect 17975 17920 18039 17924
rect 18055 17980 18119 17984
rect 18055 17924 18059 17980
rect 18059 17924 18115 17980
rect 18115 17924 18119 17980
rect 18055 17920 18119 17924
rect 18135 17980 18199 17984
rect 18135 17924 18139 17980
rect 18139 17924 18195 17980
rect 18195 17924 18199 17980
rect 18135 17920 18199 17924
rect 7729 17436 7793 17440
rect 7729 17380 7733 17436
rect 7733 17380 7789 17436
rect 7789 17380 7793 17436
rect 7729 17376 7793 17380
rect 7809 17436 7873 17440
rect 7809 17380 7813 17436
rect 7813 17380 7869 17436
rect 7869 17380 7873 17436
rect 7809 17376 7873 17380
rect 7889 17436 7953 17440
rect 7889 17380 7893 17436
rect 7893 17380 7949 17436
rect 7949 17380 7953 17436
rect 7889 17376 7953 17380
rect 7969 17436 8033 17440
rect 7969 17380 7973 17436
rect 7973 17380 8029 17436
rect 8029 17380 8033 17436
rect 7969 17376 8033 17380
rect 14506 17436 14570 17440
rect 14506 17380 14510 17436
rect 14510 17380 14566 17436
rect 14566 17380 14570 17436
rect 14506 17376 14570 17380
rect 14586 17436 14650 17440
rect 14586 17380 14590 17436
rect 14590 17380 14646 17436
rect 14646 17380 14650 17436
rect 14586 17376 14650 17380
rect 14666 17436 14730 17440
rect 14666 17380 14670 17436
rect 14670 17380 14726 17436
rect 14726 17380 14730 17436
rect 14666 17376 14730 17380
rect 14746 17436 14810 17440
rect 14746 17380 14750 17436
rect 14750 17380 14806 17436
rect 14806 17380 14810 17436
rect 14746 17376 14810 17380
rect 4340 16892 4404 16896
rect 4340 16836 4344 16892
rect 4344 16836 4400 16892
rect 4400 16836 4404 16892
rect 4340 16832 4404 16836
rect 4420 16892 4484 16896
rect 4420 16836 4424 16892
rect 4424 16836 4480 16892
rect 4480 16836 4484 16892
rect 4420 16832 4484 16836
rect 4500 16892 4564 16896
rect 4500 16836 4504 16892
rect 4504 16836 4560 16892
rect 4560 16836 4564 16892
rect 4500 16832 4564 16836
rect 4580 16892 4644 16896
rect 4580 16836 4584 16892
rect 4584 16836 4640 16892
rect 4640 16836 4644 16892
rect 4580 16832 4644 16836
rect 11118 16892 11182 16896
rect 11118 16836 11122 16892
rect 11122 16836 11178 16892
rect 11178 16836 11182 16892
rect 11118 16832 11182 16836
rect 11198 16892 11262 16896
rect 11198 16836 11202 16892
rect 11202 16836 11258 16892
rect 11258 16836 11262 16892
rect 11198 16832 11262 16836
rect 11278 16892 11342 16896
rect 11278 16836 11282 16892
rect 11282 16836 11338 16892
rect 11338 16836 11342 16892
rect 11278 16832 11342 16836
rect 11358 16892 11422 16896
rect 11358 16836 11362 16892
rect 11362 16836 11418 16892
rect 11418 16836 11422 16892
rect 11358 16832 11422 16836
rect 17895 16892 17959 16896
rect 17895 16836 17899 16892
rect 17899 16836 17955 16892
rect 17955 16836 17959 16892
rect 17895 16832 17959 16836
rect 17975 16892 18039 16896
rect 17975 16836 17979 16892
rect 17979 16836 18035 16892
rect 18035 16836 18039 16892
rect 17975 16832 18039 16836
rect 18055 16892 18119 16896
rect 18055 16836 18059 16892
rect 18059 16836 18115 16892
rect 18115 16836 18119 16892
rect 18055 16832 18119 16836
rect 18135 16892 18199 16896
rect 18135 16836 18139 16892
rect 18139 16836 18195 16892
rect 18195 16836 18199 16892
rect 18135 16832 18199 16836
rect 17724 16628 17788 16692
rect 8156 16492 8220 16556
rect 9260 16552 9324 16556
rect 9260 16496 9310 16552
rect 9310 16496 9324 16552
rect 9260 16492 9324 16496
rect 7729 16348 7793 16352
rect 7729 16292 7733 16348
rect 7733 16292 7789 16348
rect 7789 16292 7793 16348
rect 7729 16288 7793 16292
rect 7809 16348 7873 16352
rect 7809 16292 7813 16348
rect 7813 16292 7869 16348
rect 7869 16292 7873 16348
rect 7809 16288 7873 16292
rect 7889 16348 7953 16352
rect 7889 16292 7893 16348
rect 7893 16292 7949 16348
rect 7949 16292 7953 16348
rect 7889 16288 7953 16292
rect 7969 16348 8033 16352
rect 7969 16292 7973 16348
rect 7973 16292 8029 16348
rect 8029 16292 8033 16348
rect 7969 16288 8033 16292
rect 14506 16348 14570 16352
rect 14506 16292 14510 16348
rect 14510 16292 14566 16348
rect 14566 16292 14570 16348
rect 14506 16288 14570 16292
rect 14586 16348 14650 16352
rect 14586 16292 14590 16348
rect 14590 16292 14646 16348
rect 14646 16292 14650 16348
rect 14586 16288 14650 16292
rect 14666 16348 14730 16352
rect 14666 16292 14670 16348
rect 14670 16292 14726 16348
rect 14726 16292 14730 16348
rect 14666 16288 14730 16292
rect 14746 16348 14810 16352
rect 14746 16292 14750 16348
rect 14750 16292 14806 16348
rect 14806 16292 14810 16348
rect 14746 16288 14810 16292
rect 4340 15804 4404 15808
rect 4340 15748 4344 15804
rect 4344 15748 4400 15804
rect 4400 15748 4404 15804
rect 4340 15744 4404 15748
rect 4420 15804 4484 15808
rect 4420 15748 4424 15804
rect 4424 15748 4480 15804
rect 4480 15748 4484 15804
rect 4420 15744 4484 15748
rect 4500 15804 4564 15808
rect 4500 15748 4504 15804
rect 4504 15748 4560 15804
rect 4560 15748 4564 15804
rect 4500 15744 4564 15748
rect 4580 15804 4644 15808
rect 4580 15748 4584 15804
rect 4584 15748 4640 15804
rect 4640 15748 4644 15804
rect 4580 15744 4644 15748
rect 11118 15804 11182 15808
rect 11118 15748 11122 15804
rect 11122 15748 11178 15804
rect 11178 15748 11182 15804
rect 11118 15744 11182 15748
rect 11198 15804 11262 15808
rect 11198 15748 11202 15804
rect 11202 15748 11258 15804
rect 11258 15748 11262 15804
rect 11198 15744 11262 15748
rect 11278 15804 11342 15808
rect 11278 15748 11282 15804
rect 11282 15748 11338 15804
rect 11338 15748 11342 15804
rect 11278 15744 11342 15748
rect 11358 15804 11422 15808
rect 11358 15748 11362 15804
rect 11362 15748 11418 15804
rect 11418 15748 11422 15804
rect 11358 15744 11422 15748
rect 17895 15804 17959 15808
rect 17895 15748 17899 15804
rect 17899 15748 17955 15804
rect 17955 15748 17959 15804
rect 17895 15744 17959 15748
rect 17975 15804 18039 15808
rect 17975 15748 17979 15804
rect 17979 15748 18035 15804
rect 18035 15748 18039 15804
rect 17975 15744 18039 15748
rect 18055 15804 18119 15808
rect 18055 15748 18059 15804
rect 18059 15748 18115 15804
rect 18115 15748 18119 15804
rect 18055 15744 18119 15748
rect 18135 15804 18199 15808
rect 18135 15748 18139 15804
rect 18139 15748 18195 15804
rect 18195 15748 18199 15804
rect 18135 15744 18199 15748
rect 7729 15260 7793 15264
rect 7729 15204 7733 15260
rect 7733 15204 7789 15260
rect 7789 15204 7793 15260
rect 7729 15200 7793 15204
rect 7809 15260 7873 15264
rect 7809 15204 7813 15260
rect 7813 15204 7869 15260
rect 7869 15204 7873 15260
rect 7809 15200 7873 15204
rect 7889 15260 7953 15264
rect 7889 15204 7893 15260
rect 7893 15204 7949 15260
rect 7949 15204 7953 15260
rect 7889 15200 7953 15204
rect 7969 15260 8033 15264
rect 7969 15204 7973 15260
rect 7973 15204 8029 15260
rect 8029 15204 8033 15260
rect 7969 15200 8033 15204
rect 14506 15260 14570 15264
rect 14506 15204 14510 15260
rect 14510 15204 14566 15260
rect 14566 15204 14570 15260
rect 14506 15200 14570 15204
rect 14586 15260 14650 15264
rect 14586 15204 14590 15260
rect 14590 15204 14646 15260
rect 14646 15204 14650 15260
rect 14586 15200 14650 15204
rect 14666 15260 14730 15264
rect 14666 15204 14670 15260
rect 14670 15204 14726 15260
rect 14726 15204 14730 15260
rect 14666 15200 14730 15204
rect 14746 15260 14810 15264
rect 14746 15204 14750 15260
rect 14750 15204 14806 15260
rect 14806 15204 14810 15260
rect 14746 15200 14810 15204
rect 4340 14716 4404 14720
rect 4340 14660 4344 14716
rect 4344 14660 4400 14716
rect 4400 14660 4404 14716
rect 4340 14656 4404 14660
rect 4420 14716 4484 14720
rect 4420 14660 4424 14716
rect 4424 14660 4480 14716
rect 4480 14660 4484 14716
rect 4420 14656 4484 14660
rect 4500 14716 4564 14720
rect 4500 14660 4504 14716
rect 4504 14660 4560 14716
rect 4560 14660 4564 14716
rect 4500 14656 4564 14660
rect 4580 14716 4644 14720
rect 4580 14660 4584 14716
rect 4584 14660 4640 14716
rect 4640 14660 4644 14716
rect 4580 14656 4644 14660
rect 11118 14716 11182 14720
rect 11118 14660 11122 14716
rect 11122 14660 11178 14716
rect 11178 14660 11182 14716
rect 11118 14656 11182 14660
rect 11198 14716 11262 14720
rect 11198 14660 11202 14716
rect 11202 14660 11258 14716
rect 11258 14660 11262 14716
rect 11198 14656 11262 14660
rect 11278 14716 11342 14720
rect 11278 14660 11282 14716
rect 11282 14660 11338 14716
rect 11338 14660 11342 14716
rect 11278 14656 11342 14660
rect 11358 14716 11422 14720
rect 11358 14660 11362 14716
rect 11362 14660 11418 14716
rect 11418 14660 11422 14716
rect 11358 14656 11422 14660
rect 17895 14716 17959 14720
rect 17895 14660 17899 14716
rect 17899 14660 17955 14716
rect 17955 14660 17959 14716
rect 17895 14656 17959 14660
rect 17975 14716 18039 14720
rect 17975 14660 17979 14716
rect 17979 14660 18035 14716
rect 18035 14660 18039 14716
rect 17975 14656 18039 14660
rect 18055 14716 18119 14720
rect 18055 14660 18059 14716
rect 18059 14660 18115 14716
rect 18115 14660 18119 14716
rect 18055 14656 18119 14660
rect 18135 14716 18199 14720
rect 18135 14660 18139 14716
rect 18139 14660 18195 14716
rect 18195 14660 18199 14716
rect 18135 14656 18199 14660
rect 7729 14172 7793 14176
rect 7729 14116 7733 14172
rect 7733 14116 7789 14172
rect 7789 14116 7793 14172
rect 7729 14112 7793 14116
rect 7809 14172 7873 14176
rect 7809 14116 7813 14172
rect 7813 14116 7869 14172
rect 7869 14116 7873 14172
rect 7809 14112 7873 14116
rect 7889 14172 7953 14176
rect 7889 14116 7893 14172
rect 7893 14116 7949 14172
rect 7949 14116 7953 14172
rect 7889 14112 7953 14116
rect 7969 14172 8033 14176
rect 7969 14116 7973 14172
rect 7973 14116 8029 14172
rect 8029 14116 8033 14172
rect 7969 14112 8033 14116
rect 14506 14172 14570 14176
rect 14506 14116 14510 14172
rect 14510 14116 14566 14172
rect 14566 14116 14570 14172
rect 14506 14112 14570 14116
rect 14586 14172 14650 14176
rect 14586 14116 14590 14172
rect 14590 14116 14646 14172
rect 14646 14116 14650 14172
rect 14586 14112 14650 14116
rect 14666 14172 14730 14176
rect 14666 14116 14670 14172
rect 14670 14116 14726 14172
rect 14726 14116 14730 14172
rect 14666 14112 14730 14116
rect 14746 14172 14810 14176
rect 14746 14116 14750 14172
rect 14750 14116 14806 14172
rect 14806 14116 14810 14172
rect 14746 14112 14810 14116
rect 9260 14104 9324 14108
rect 9260 14048 9274 14104
rect 9274 14048 9324 14104
rect 9260 14044 9324 14048
rect 17724 13908 17788 13972
rect 4340 13628 4404 13632
rect 4340 13572 4344 13628
rect 4344 13572 4400 13628
rect 4400 13572 4404 13628
rect 4340 13568 4404 13572
rect 4420 13628 4484 13632
rect 4420 13572 4424 13628
rect 4424 13572 4480 13628
rect 4480 13572 4484 13628
rect 4420 13568 4484 13572
rect 4500 13628 4564 13632
rect 4500 13572 4504 13628
rect 4504 13572 4560 13628
rect 4560 13572 4564 13628
rect 4500 13568 4564 13572
rect 4580 13628 4644 13632
rect 4580 13572 4584 13628
rect 4584 13572 4640 13628
rect 4640 13572 4644 13628
rect 4580 13568 4644 13572
rect 11118 13628 11182 13632
rect 11118 13572 11122 13628
rect 11122 13572 11178 13628
rect 11178 13572 11182 13628
rect 11118 13568 11182 13572
rect 11198 13628 11262 13632
rect 11198 13572 11202 13628
rect 11202 13572 11258 13628
rect 11258 13572 11262 13628
rect 11198 13568 11262 13572
rect 11278 13628 11342 13632
rect 11278 13572 11282 13628
rect 11282 13572 11338 13628
rect 11338 13572 11342 13628
rect 11278 13568 11342 13572
rect 11358 13628 11422 13632
rect 11358 13572 11362 13628
rect 11362 13572 11418 13628
rect 11418 13572 11422 13628
rect 11358 13568 11422 13572
rect 17895 13628 17959 13632
rect 17895 13572 17899 13628
rect 17899 13572 17955 13628
rect 17955 13572 17959 13628
rect 17895 13568 17959 13572
rect 17975 13628 18039 13632
rect 17975 13572 17979 13628
rect 17979 13572 18035 13628
rect 18035 13572 18039 13628
rect 17975 13568 18039 13572
rect 18055 13628 18119 13632
rect 18055 13572 18059 13628
rect 18059 13572 18115 13628
rect 18115 13572 18119 13628
rect 18055 13568 18119 13572
rect 18135 13628 18199 13632
rect 18135 13572 18139 13628
rect 18139 13572 18195 13628
rect 18195 13572 18199 13628
rect 18135 13568 18199 13572
rect 14964 13364 15028 13428
rect 7729 13084 7793 13088
rect 7729 13028 7733 13084
rect 7733 13028 7789 13084
rect 7789 13028 7793 13084
rect 7729 13024 7793 13028
rect 7809 13084 7873 13088
rect 7809 13028 7813 13084
rect 7813 13028 7869 13084
rect 7869 13028 7873 13084
rect 7809 13024 7873 13028
rect 7889 13084 7953 13088
rect 7889 13028 7893 13084
rect 7893 13028 7949 13084
rect 7949 13028 7953 13084
rect 7889 13024 7953 13028
rect 7969 13084 8033 13088
rect 7969 13028 7973 13084
rect 7973 13028 8029 13084
rect 8029 13028 8033 13084
rect 7969 13024 8033 13028
rect 14506 13084 14570 13088
rect 14506 13028 14510 13084
rect 14510 13028 14566 13084
rect 14566 13028 14570 13084
rect 14506 13024 14570 13028
rect 14586 13084 14650 13088
rect 14586 13028 14590 13084
rect 14590 13028 14646 13084
rect 14646 13028 14650 13084
rect 14586 13024 14650 13028
rect 14666 13084 14730 13088
rect 14666 13028 14670 13084
rect 14670 13028 14726 13084
rect 14726 13028 14730 13084
rect 14666 13024 14730 13028
rect 14746 13084 14810 13088
rect 14746 13028 14750 13084
rect 14750 13028 14806 13084
rect 14806 13028 14810 13084
rect 14746 13024 14810 13028
rect 4340 12540 4404 12544
rect 4340 12484 4344 12540
rect 4344 12484 4400 12540
rect 4400 12484 4404 12540
rect 4340 12480 4404 12484
rect 4420 12540 4484 12544
rect 4420 12484 4424 12540
rect 4424 12484 4480 12540
rect 4480 12484 4484 12540
rect 4420 12480 4484 12484
rect 4500 12540 4564 12544
rect 4500 12484 4504 12540
rect 4504 12484 4560 12540
rect 4560 12484 4564 12540
rect 4500 12480 4564 12484
rect 4580 12540 4644 12544
rect 4580 12484 4584 12540
rect 4584 12484 4640 12540
rect 4640 12484 4644 12540
rect 4580 12480 4644 12484
rect 11118 12540 11182 12544
rect 11118 12484 11122 12540
rect 11122 12484 11178 12540
rect 11178 12484 11182 12540
rect 11118 12480 11182 12484
rect 11198 12540 11262 12544
rect 11198 12484 11202 12540
rect 11202 12484 11258 12540
rect 11258 12484 11262 12540
rect 11198 12480 11262 12484
rect 11278 12540 11342 12544
rect 11278 12484 11282 12540
rect 11282 12484 11338 12540
rect 11338 12484 11342 12540
rect 11278 12480 11342 12484
rect 11358 12540 11422 12544
rect 11358 12484 11362 12540
rect 11362 12484 11418 12540
rect 11418 12484 11422 12540
rect 11358 12480 11422 12484
rect 17895 12540 17959 12544
rect 17895 12484 17899 12540
rect 17899 12484 17955 12540
rect 17955 12484 17959 12540
rect 17895 12480 17959 12484
rect 17975 12540 18039 12544
rect 17975 12484 17979 12540
rect 17979 12484 18035 12540
rect 18035 12484 18039 12540
rect 17975 12480 18039 12484
rect 18055 12540 18119 12544
rect 18055 12484 18059 12540
rect 18059 12484 18115 12540
rect 18115 12484 18119 12540
rect 18055 12480 18119 12484
rect 18135 12540 18199 12544
rect 18135 12484 18139 12540
rect 18139 12484 18195 12540
rect 18195 12484 18199 12540
rect 18135 12480 18199 12484
rect 8156 12412 8220 12476
rect 7729 11996 7793 12000
rect 7729 11940 7733 11996
rect 7733 11940 7789 11996
rect 7789 11940 7793 11996
rect 7729 11936 7793 11940
rect 7809 11996 7873 12000
rect 7809 11940 7813 11996
rect 7813 11940 7869 11996
rect 7869 11940 7873 11996
rect 7809 11936 7873 11940
rect 7889 11996 7953 12000
rect 7889 11940 7893 11996
rect 7893 11940 7949 11996
rect 7949 11940 7953 11996
rect 7889 11936 7953 11940
rect 7969 11996 8033 12000
rect 7969 11940 7973 11996
rect 7973 11940 8029 11996
rect 8029 11940 8033 11996
rect 7969 11936 8033 11940
rect 14506 11996 14570 12000
rect 14506 11940 14510 11996
rect 14510 11940 14566 11996
rect 14566 11940 14570 11996
rect 14506 11936 14570 11940
rect 14586 11996 14650 12000
rect 14586 11940 14590 11996
rect 14590 11940 14646 11996
rect 14646 11940 14650 11996
rect 14586 11936 14650 11940
rect 14666 11996 14730 12000
rect 14666 11940 14670 11996
rect 14670 11940 14726 11996
rect 14726 11940 14730 11996
rect 14666 11936 14730 11940
rect 14746 11996 14810 12000
rect 14746 11940 14750 11996
rect 14750 11940 14806 11996
rect 14806 11940 14810 11996
rect 14746 11936 14810 11940
rect 4340 11452 4404 11456
rect 4340 11396 4344 11452
rect 4344 11396 4400 11452
rect 4400 11396 4404 11452
rect 4340 11392 4404 11396
rect 4420 11452 4484 11456
rect 4420 11396 4424 11452
rect 4424 11396 4480 11452
rect 4480 11396 4484 11452
rect 4420 11392 4484 11396
rect 4500 11452 4564 11456
rect 4500 11396 4504 11452
rect 4504 11396 4560 11452
rect 4560 11396 4564 11452
rect 4500 11392 4564 11396
rect 4580 11452 4644 11456
rect 4580 11396 4584 11452
rect 4584 11396 4640 11452
rect 4640 11396 4644 11452
rect 4580 11392 4644 11396
rect 11118 11452 11182 11456
rect 11118 11396 11122 11452
rect 11122 11396 11178 11452
rect 11178 11396 11182 11452
rect 11118 11392 11182 11396
rect 11198 11452 11262 11456
rect 11198 11396 11202 11452
rect 11202 11396 11258 11452
rect 11258 11396 11262 11452
rect 11198 11392 11262 11396
rect 11278 11452 11342 11456
rect 11278 11396 11282 11452
rect 11282 11396 11338 11452
rect 11338 11396 11342 11452
rect 11278 11392 11342 11396
rect 11358 11452 11422 11456
rect 11358 11396 11362 11452
rect 11362 11396 11418 11452
rect 11418 11396 11422 11452
rect 11358 11392 11422 11396
rect 17895 11452 17959 11456
rect 17895 11396 17899 11452
rect 17899 11396 17955 11452
rect 17955 11396 17959 11452
rect 17895 11392 17959 11396
rect 17975 11452 18039 11456
rect 17975 11396 17979 11452
rect 17979 11396 18035 11452
rect 18035 11396 18039 11452
rect 17975 11392 18039 11396
rect 18055 11452 18119 11456
rect 18055 11396 18059 11452
rect 18059 11396 18115 11452
rect 18115 11396 18119 11452
rect 18055 11392 18119 11396
rect 18135 11452 18199 11456
rect 18135 11396 18139 11452
rect 18139 11396 18195 11452
rect 18195 11396 18199 11452
rect 18135 11392 18199 11396
rect 7729 10908 7793 10912
rect 7729 10852 7733 10908
rect 7733 10852 7789 10908
rect 7789 10852 7793 10908
rect 7729 10848 7793 10852
rect 7809 10908 7873 10912
rect 7809 10852 7813 10908
rect 7813 10852 7869 10908
rect 7869 10852 7873 10908
rect 7809 10848 7873 10852
rect 7889 10908 7953 10912
rect 7889 10852 7893 10908
rect 7893 10852 7949 10908
rect 7949 10852 7953 10908
rect 7889 10848 7953 10852
rect 7969 10908 8033 10912
rect 7969 10852 7973 10908
rect 7973 10852 8029 10908
rect 8029 10852 8033 10908
rect 7969 10848 8033 10852
rect 14506 10908 14570 10912
rect 14506 10852 14510 10908
rect 14510 10852 14566 10908
rect 14566 10852 14570 10908
rect 14506 10848 14570 10852
rect 14586 10908 14650 10912
rect 14586 10852 14590 10908
rect 14590 10852 14646 10908
rect 14646 10852 14650 10908
rect 14586 10848 14650 10852
rect 14666 10908 14730 10912
rect 14666 10852 14670 10908
rect 14670 10852 14726 10908
rect 14726 10852 14730 10908
rect 14666 10848 14730 10852
rect 14746 10908 14810 10912
rect 14746 10852 14750 10908
rect 14750 10852 14806 10908
rect 14806 10852 14810 10908
rect 14746 10848 14810 10852
rect 4340 10364 4404 10368
rect 4340 10308 4344 10364
rect 4344 10308 4400 10364
rect 4400 10308 4404 10364
rect 4340 10304 4404 10308
rect 4420 10364 4484 10368
rect 4420 10308 4424 10364
rect 4424 10308 4480 10364
rect 4480 10308 4484 10364
rect 4420 10304 4484 10308
rect 4500 10364 4564 10368
rect 4500 10308 4504 10364
rect 4504 10308 4560 10364
rect 4560 10308 4564 10364
rect 4500 10304 4564 10308
rect 4580 10364 4644 10368
rect 4580 10308 4584 10364
rect 4584 10308 4640 10364
rect 4640 10308 4644 10364
rect 4580 10304 4644 10308
rect 11118 10364 11182 10368
rect 11118 10308 11122 10364
rect 11122 10308 11178 10364
rect 11178 10308 11182 10364
rect 11118 10304 11182 10308
rect 11198 10364 11262 10368
rect 11198 10308 11202 10364
rect 11202 10308 11258 10364
rect 11258 10308 11262 10364
rect 11198 10304 11262 10308
rect 11278 10364 11342 10368
rect 11278 10308 11282 10364
rect 11282 10308 11338 10364
rect 11338 10308 11342 10364
rect 11278 10304 11342 10308
rect 11358 10364 11422 10368
rect 11358 10308 11362 10364
rect 11362 10308 11418 10364
rect 11418 10308 11422 10364
rect 11358 10304 11422 10308
rect 17895 10364 17959 10368
rect 17895 10308 17899 10364
rect 17899 10308 17955 10364
rect 17955 10308 17959 10364
rect 17895 10304 17959 10308
rect 17975 10364 18039 10368
rect 17975 10308 17979 10364
rect 17979 10308 18035 10364
rect 18035 10308 18039 10364
rect 17975 10304 18039 10308
rect 18055 10364 18119 10368
rect 18055 10308 18059 10364
rect 18059 10308 18115 10364
rect 18115 10308 18119 10364
rect 18055 10304 18119 10308
rect 18135 10364 18199 10368
rect 18135 10308 18139 10364
rect 18139 10308 18195 10364
rect 18195 10308 18199 10364
rect 18135 10304 18199 10308
rect 7729 9820 7793 9824
rect 7729 9764 7733 9820
rect 7733 9764 7789 9820
rect 7789 9764 7793 9820
rect 7729 9760 7793 9764
rect 7809 9820 7873 9824
rect 7809 9764 7813 9820
rect 7813 9764 7869 9820
rect 7869 9764 7873 9820
rect 7809 9760 7873 9764
rect 7889 9820 7953 9824
rect 7889 9764 7893 9820
rect 7893 9764 7949 9820
rect 7949 9764 7953 9820
rect 7889 9760 7953 9764
rect 7969 9820 8033 9824
rect 7969 9764 7973 9820
rect 7973 9764 8029 9820
rect 8029 9764 8033 9820
rect 7969 9760 8033 9764
rect 14506 9820 14570 9824
rect 14506 9764 14510 9820
rect 14510 9764 14566 9820
rect 14566 9764 14570 9820
rect 14506 9760 14570 9764
rect 14586 9820 14650 9824
rect 14586 9764 14590 9820
rect 14590 9764 14646 9820
rect 14646 9764 14650 9820
rect 14586 9760 14650 9764
rect 14666 9820 14730 9824
rect 14666 9764 14670 9820
rect 14670 9764 14726 9820
rect 14726 9764 14730 9820
rect 14666 9760 14730 9764
rect 14746 9820 14810 9824
rect 14746 9764 14750 9820
rect 14750 9764 14806 9820
rect 14806 9764 14810 9820
rect 14746 9760 14810 9764
rect 20300 9420 20364 9484
rect 4340 9276 4404 9280
rect 4340 9220 4344 9276
rect 4344 9220 4400 9276
rect 4400 9220 4404 9276
rect 4340 9216 4404 9220
rect 4420 9276 4484 9280
rect 4420 9220 4424 9276
rect 4424 9220 4480 9276
rect 4480 9220 4484 9276
rect 4420 9216 4484 9220
rect 4500 9276 4564 9280
rect 4500 9220 4504 9276
rect 4504 9220 4560 9276
rect 4560 9220 4564 9276
rect 4500 9216 4564 9220
rect 4580 9276 4644 9280
rect 4580 9220 4584 9276
rect 4584 9220 4640 9276
rect 4640 9220 4644 9276
rect 4580 9216 4644 9220
rect 11118 9276 11182 9280
rect 11118 9220 11122 9276
rect 11122 9220 11178 9276
rect 11178 9220 11182 9276
rect 11118 9216 11182 9220
rect 11198 9276 11262 9280
rect 11198 9220 11202 9276
rect 11202 9220 11258 9276
rect 11258 9220 11262 9276
rect 11198 9216 11262 9220
rect 11278 9276 11342 9280
rect 11278 9220 11282 9276
rect 11282 9220 11338 9276
rect 11338 9220 11342 9276
rect 11278 9216 11342 9220
rect 11358 9276 11422 9280
rect 11358 9220 11362 9276
rect 11362 9220 11418 9276
rect 11418 9220 11422 9276
rect 11358 9216 11422 9220
rect 17895 9276 17959 9280
rect 17895 9220 17899 9276
rect 17899 9220 17955 9276
rect 17955 9220 17959 9276
rect 17895 9216 17959 9220
rect 17975 9276 18039 9280
rect 17975 9220 17979 9276
rect 17979 9220 18035 9276
rect 18035 9220 18039 9276
rect 17975 9216 18039 9220
rect 18055 9276 18119 9280
rect 18055 9220 18059 9276
rect 18059 9220 18115 9276
rect 18115 9220 18119 9276
rect 18055 9216 18119 9220
rect 18135 9276 18199 9280
rect 18135 9220 18139 9276
rect 18139 9220 18195 9276
rect 18195 9220 18199 9276
rect 18135 9216 18199 9220
rect 19932 9012 19996 9076
rect 7729 8732 7793 8736
rect 7729 8676 7733 8732
rect 7733 8676 7789 8732
rect 7789 8676 7793 8732
rect 7729 8672 7793 8676
rect 7809 8732 7873 8736
rect 7809 8676 7813 8732
rect 7813 8676 7869 8732
rect 7869 8676 7873 8732
rect 7809 8672 7873 8676
rect 7889 8732 7953 8736
rect 7889 8676 7893 8732
rect 7893 8676 7949 8732
rect 7949 8676 7953 8732
rect 7889 8672 7953 8676
rect 7969 8732 8033 8736
rect 7969 8676 7973 8732
rect 7973 8676 8029 8732
rect 8029 8676 8033 8732
rect 7969 8672 8033 8676
rect 14506 8732 14570 8736
rect 14506 8676 14510 8732
rect 14510 8676 14566 8732
rect 14566 8676 14570 8732
rect 14506 8672 14570 8676
rect 14586 8732 14650 8736
rect 14586 8676 14590 8732
rect 14590 8676 14646 8732
rect 14646 8676 14650 8732
rect 14586 8672 14650 8676
rect 14666 8732 14730 8736
rect 14666 8676 14670 8732
rect 14670 8676 14726 8732
rect 14726 8676 14730 8732
rect 14666 8672 14730 8676
rect 14746 8732 14810 8736
rect 14746 8676 14750 8732
rect 14750 8676 14806 8732
rect 14806 8676 14810 8732
rect 14746 8672 14810 8676
rect 4340 8188 4404 8192
rect 4340 8132 4344 8188
rect 4344 8132 4400 8188
rect 4400 8132 4404 8188
rect 4340 8128 4404 8132
rect 4420 8188 4484 8192
rect 4420 8132 4424 8188
rect 4424 8132 4480 8188
rect 4480 8132 4484 8188
rect 4420 8128 4484 8132
rect 4500 8188 4564 8192
rect 4500 8132 4504 8188
rect 4504 8132 4560 8188
rect 4560 8132 4564 8188
rect 4500 8128 4564 8132
rect 4580 8188 4644 8192
rect 4580 8132 4584 8188
rect 4584 8132 4640 8188
rect 4640 8132 4644 8188
rect 4580 8128 4644 8132
rect 11118 8188 11182 8192
rect 11118 8132 11122 8188
rect 11122 8132 11178 8188
rect 11178 8132 11182 8188
rect 11118 8128 11182 8132
rect 11198 8188 11262 8192
rect 11198 8132 11202 8188
rect 11202 8132 11258 8188
rect 11258 8132 11262 8188
rect 11198 8128 11262 8132
rect 11278 8188 11342 8192
rect 11278 8132 11282 8188
rect 11282 8132 11338 8188
rect 11338 8132 11342 8188
rect 11278 8128 11342 8132
rect 11358 8188 11422 8192
rect 11358 8132 11362 8188
rect 11362 8132 11418 8188
rect 11418 8132 11422 8188
rect 11358 8128 11422 8132
rect 17895 8188 17959 8192
rect 17895 8132 17899 8188
rect 17899 8132 17955 8188
rect 17955 8132 17959 8188
rect 17895 8128 17959 8132
rect 17975 8188 18039 8192
rect 17975 8132 17979 8188
rect 17979 8132 18035 8188
rect 18035 8132 18039 8188
rect 17975 8128 18039 8132
rect 18055 8188 18119 8192
rect 18055 8132 18059 8188
rect 18059 8132 18115 8188
rect 18115 8132 18119 8188
rect 18055 8128 18119 8132
rect 18135 8188 18199 8192
rect 18135 8132 18139 8188
rect 18139 8132 18195 8188
rect 18195 8132 18199 8188
rect 18135 8128 18199 8132
rect 7729 7644 7793 7648
rect 7729 7588 7733 7644
rect 7733 7588 7789 7644
rect 7789 7588 7793 7644
rect 7729 7584 7793 7588
rect 7809 7644 7873 7648
rect 7809 7588 7813 7644
rect 7813 7588 7869 7644
rect 7869 7588 7873 7644
rect 7809 7584 7873 7588
rect 7889 7644 7953 7648
rect 7889 7588 7893 7644
rect 7893 7588 7949 7644
rect 7949 7588 7953 7644
rect 7889 7584 7953 7588
rect 7969 7644 8033 7648
rect 7969 7588 7973 7644
rect 7973 7588 8029 7644
rect 8029 7588 8033 7644
rect 7969 7584 8033 7588
rect 14506 7644 14570 7648
rect 14506 7588 14510 7644
rect 14510 7588 14566 7644
rect 14566 7588 14570 7644
rect 14506 7584 14570 7588
rect 14586 7644 14650 7648
rect 14586 7588 14590 7644
rect 14590 7588 14646 7644
rect 14646 7588 14650 7644
rect 14586 7584 14650 7588
rect 14666 7644 14730 7648
rect 14666 7588 14670 7644
rect 14670 7588 14726 7644
rect 14726 7588 14730 7644
rect 14666 7584 14730 7588
rect 14746 7644 14810 7648
rect 14746 7588 14750 7644
rect 14750 7588 14806 7644
rect 14806 7588 14810 7644
rect 14746 7584 14810 7588
rect 20484 7380 20548 7444
rect 4340 7100 4404 7104
rect 4340 7044 4344 7100
rect 4344 7044 4400 7100
rect 4400 7044 4404 7100
rect 4340 7040 4404 7044
rect 4420 7100 4484 7104
rect 4420 7044 4424 7100
rect 4424 7044 4480 7100
rect 4480 7044 4484 7100
rect 4420 7040 4484 7044
rect 4500 7100 4564 7104
rect 4500 7044 4504 7100
rect 4504 7044 4560 7100
rect 4560 7044 4564 7100
rect 4500 7040 4564 7044
rect 4580 7100 4644 7104
rect 4580 7044 4584 7100
rect 4584 7044 4640 7100
rect 4640 7044 4644 7100
rect 4580 7040 4644 7044
rect 11118 7100 11182 7104
rect 11118 7044 11122 7100
rect 11122 7044 11178 7100
rect 11178 7044 11182 7100
rect 11118 7040 11182 7044
rect 11198 7100 11262 7104
rect 11198 7044 11202 7100
rect 11202 7044 11258 7100
rect 11258 7044 11262 7100
rect 11198 7040 11262 7044
rect 11278 7100 11342 7104
rect 11278 7044 11282 7100
rect 11282 7044 11338 7100
rect 11338 7044 11342 7100
rect 11278 7040 11342 7044
rect 11358 7100 11422 7104
rect 11358 7044 11362 7100
rect 11362 7044 11418 7100
rect 11418 7044 11422 7100
rect 11358 7040 11422 7044
rect 17895 7100 17959 7104
rect 17895 7044 17899 7100
rect 17899 7044 17955 7100
rect 17955 7044 17959 7100
rect 17895 7040 17959 7044
rect 17975 7100 18039 7104
rect 17975 7044 17979 7100
rect 17979 7044 18035 7100
rect 18035 7044 18039 7100
rect 17975 7040 18039 7044
rect 18055 7100 18119 7104
rect 18055 7044 18059 7100
rect 18059 7044 18115 7100
rect 18115 7044 18119 7100
rect 18055 7040 18119 7044
rect 18135 7100 18199 7104
rect 18135 7044 18139 7100
rect 18139 7044 18195 7100
rect 18195 7044 18199 7100
rect 18135 7040 18199 7044
rect 8156 6972 8220 7036
rect 7729 6556 7793 6560
rect 7729 6500 7733 6556
rect 7733 6500 7789 6556
rect 7789 6500 7793 6556
rect 7729 6496 7793 6500
rect 7809 6556 7873 6560
rect 7809 6500 7813 6556
rect 7813 6500 7869 6556
rect 7869 6500 7873 6556
rect 7809 6496 7873 6500
rect 7889 6556 7953 6560
rect 7889 6500 7893 6556
rect 7893 6500 7949 6556
rect 7949 6500 7953 6556
rect 7889 6496 7953 6500
rect 7969 6556 8033 6560
rect 7969 6500 7973 6556
rect 7973 6500 8029 6556
rect 8029 6500 8033 6556
rect 7969 6496 8033 6500
rect 14506 6556 14570 6560
rect 14506 6500 14510 6556
rect 14510 6500 14566 6556
rect 14566 6500 14570 6556
rect 14506 6496 14570 6500
rect 14586 6556 14650 6560
rect 14586 6500 14590 6556
rect 14590 6500 14646 6556
rect 14646 6500 14650 6556
rect 14586 6496 14650 6500
rect 14666 6556 14730 6560
rect 14666 6500 14670 6556
rect 14670 6500 14726 6556
rect 14726 6500 14730 6556
rect 14666 6496 14730 6500
rect 14746 6556 14810 6560
rect 14746 6500 14750 6556
rect 14750 6500 14806 6556
rect 14806 6500 14810 6556
rect 14746 6496 14810 6500
rect 4340 6012 4404 6016
rect 4340 5956 4344 6012
rect 4344 5956 4400 6012
rect 4400 5956 4404 6012
rect 4340 5952 4404 5956
rect 4420 6012 4484 6016
rect 4420 5956 4424 6012
rect 4424 5956 4480 6012
rect 4480 5956 4484 6012
rect 4420 5952 4484 5956
rect 4500 6012 4564 6016
rect 4500 5956 4504 6012
rect 4504 5956 4560 6012
rect 4560 5956 4564 6012
rect 4500 5952 4564 5956
rect 4580 6012 4644 6016
rect 4580 5956 4584 6012
rect 4584 5956 4640 6012
rect 4640 5956 4644 6012
rect 4580 5952 4644 5956
rect 11118 6012 11182 6016
rect 11118 5956 11122 6012
rect 11122 5956 11178 6012
rect 11178 5956 11182 6012
rect 11118 5952 11182 5956
rect 11198 6012 11262 6016
rect 11198 5956 11202 6012
rect 11202 5956 11258 6012
rect 11258 5956 11262 6012
rect 11198 5952 11262 5956
rect 11278 6012 11342 6016
rect 11278 5956 11282 6012
rect 11282 5956 11338 6012
rect 11338 5956 11342 6012
rect 11278 5952 11342 5956
rect 11358 6012 11422 6016
rect 11358 5956 11362 6012
rect 11362 5956 11418 6012
rect 11418 5956 11422 6012
rect 11358 5952 11422 5956
rect 17895 6012 17959 6016
rect 17895 5956 17899 6012
rect 17899 5956 17955 6012
rect 17955 5956 17959 6012
rect 17895 5952 17959 5956
rect 17975 6012 18039 6016
rect 17975 5956 17979 6012
rect 17979 5956 18035 6012
rect 18035 5956 18039 6012
rect 17975 5952 18039 5956
rect 18055 6012 18119 6016
rect 18055 5956 18059 6012
rect 18059 5956 18115 6012
rect 18115 5956 18119 6012
rect 18055 5952 18119 5956
rect 18135 6012 18199 6016
rect 18135 5956 18139 6012
rect 18139 5956 18195 6012
rect 18195 5956 18199 6012
rect 18135 5952 18199 5956
rect 20116 5884 20180 5948
rect 7729 5468 7793 5472
rect 7729 5412 7733 5468
rect 7733 5412 7789 5468
rect 7789 5412 7793 5468
rect 7729 5408 7793 5412
rect 7809 5468 7873 5472
rect 7809 5412 7813 5468
rect 7813 5412 7869 5468
rect 7869 5412 7873 5468
rect 7809 5408 7873 5412
rect 7889 5468 7953 5472
rect 7889 5412 7893 5468
rect 7893 5412 7949 5468
rect 7949 5412 7953 5468
rect 7889 5408 7953 5412
rect 7969 5468 8033 5472
rect 7969 5412 7973 5468
rect 7973 5412 8029 5468
rect 8029 5412 8033 5468
rect 7969 5408 8033 5412
rect 14506 5468 14570 5472
rect 14506 5412 14510 5468
rect 14510 5412 14566 5468
rect 14566 5412 14570 5468
rect 14506 5408 14570 5412
rect 14586 5468 14650 5472
rect 14586 5412 14590 5468
rect 14590 5412 14646 5468
rect 14646 5412 14650 5468
rect 14586 5408 14650 5412
rect 14666 5468 14730 5472
rect 14666 5412 14670 5468
rect 14670 5412 14726 5468
rect 14726 5412 14730 5468
rect 14666 5408 14730 5412
rect 14746 5468 14810 5472
rect 14746 5412 14750 5468
rect 14750 5412 14806 5468
rect 14806 5412 14810 5468
rect 14746 5408 14810 5412
rect 9444 5340 9508 5404
rect 4340 4924 4404 4928
rect 4340 4868 4344 4924
rect 4344 4868 4400 4924
rect 4400 4868 4404 4924
rect 4340 4864 4404 4868
rect 4420 4924 4484 4928
rect 4420 4868 4424 4924
rect 4424 4868 4480 4924
rect 4480 4868 4484 4924
rect 4420 4864 4484 4868
rect 4500 4924 4564 4928
rect 4500 4868 4504 4924
rect 4504 4868 4560 4924
rect 4560 4868 4564 4924
rect 4500 4864 4564 4868
rect 4580 4924 4644 4928
rect 4580 4868 4584 4924
rect 4584 4868 4640 4924
rect 4640 4868 4644 4924
rect 4580 4864 4644 4868
rect 11118 4924 11182 4928
rect 11118 4868 11122 4924
rect 11122 4868 11178 4924
rect 11178 4868 11182 4924
rect 11118 4864 11182 4868
rect 11198 4924 11262 4928
rect 11198 4868 11202 4924
rect 11202 4868 11258 4924
rect 11258 4868 11262 4924
rect 11198 4864 11262 4868
rect 11278 4924 11342 4928
rect 11278 4868 11282 4924
rect 11282 4868 11338 4924
rect 11338 4868 11342 4924
rect 11278 4864 11342 4868
rect 11358 4924 11422 4928
rect 11358 4868 11362 4924
rect 11362 4868 11418 4924
rect 11418 4868 11422 4924
rect 11358 4864 11422 4868
rect 17895 4924 17959 4928
rect 17895 4868 17899 4924
rect 17899 4868 17955 4924
rect 17955 4868 17959 4924
rect 17895 4864 17959 4868
rect 17975 4924 18039 4928
rect 17975 4868 17979 4924
rect 17979 4868 18035 4924
rect 18035 4868 18039 4924
rect 17975 4864 18039 4868
rect 18055 4924 18119 4928
rect 18055 4868 18059 4924
rect 18059 4868 18115 4924
rect 18115 4868 18119 4924
rect 18055 4864 18119 4868
rect 18135 4924 18199 4928
rect 18135 4868 18139 4924
rect 18139 4868 18195 4924
rect 18195 4868 18199 4924
rect 18135 4864 18199 4868
rect 9444 4796 9508 4860
rect 7729 4380 7793 4384
rect 7729 4324 7733 4380
rect 7733 4324 7789 4380
rect 7789 4324 7793 4380
rect 7729 4320 7793 4324
rect 7809 4380 7873 4384
rect 7809 4324 7813 4380
rect 7813 4324 7869 4380
rect 7869 4324 7873 4380
rect 7809 4320 7873 4324
rect 7889 4380 7953 4384
rect 7889 4324 7893 4380
rect 7893 4324 7949 4380
rect 7949 4324 7953 4380
rect 7889 4320 7953 4324
rect 7969 4380 8033 4384
rect 7969 4324 7973 4380
rect 7973 4324 8029 4380
rect 8029 4324 8033 4380
rect 7969 4320 8033 4324
rect 14506 4380 14570 4384
rect 14506 4324 14510 4380
rect 14510 4324 14566 4380
rect 14566 4324 14570 4380
rect 14506 4320 14570 4324
rect 14586 4380 14650 4384
rect 14586 4324 14590 4380
rect 14590 4324 14646 4380
rect 14646 4324 14650 4380
rect 14586 4320 14650 4324
rect 14666 4380 14730 4384
rect 14666 4324 14670 4380
rect 14670 4324 14726 4380
rect 14726 4324 14730 4380
rect 14666 4320 14730 4324
rect 14746 4380 14810 4384
rect 14746 4324 14750 4380
rect 14750 4324 14806 4380
rect 14806 4324 14810 4380
rect 14746 4320 14810 4324
rect 4340 3836 4404 3840
rect 4340 3780 4344 3836
rect 4344 3780 4400 3836
rect 4400 3780 4404 3836
rect 4340 3776 4404 3780
rect 4420 3836 4484 3840
rect 4420 3780 4424 3836
rect 4424 3780 4480 3836
rect 4480 3780 4484 3836
rect 4420 3776 4484 3780
rect 4500 3836 4564 3840
rect 4500 3780 4504 3836
rect 4504 3780 4560 3836
rect 4560 3780 4564 3836
rect 4500 3776 4564 3780
rect 4580 3836 4644 3840
rect 4580 3780 4584 3836
rect 4584 3780 4640 3836
rect 4640 3780 4644 3836
rect 4580 3776 4644 3780
rect 11118 3836 11182 3840
rect 11118 3780 11122 3836
rect 11122 3780 11178 3836
rect 11178 3780 11182 3836
rect 11118 3776 11182 3780
rect 11198 3836 11262 3840
rect 11198 3780 11202 3836
rect 11202 3780 11258 3836
rect 11258 3780 11262 3836
rect 11198 3776 11262 3780
rect 11278 3836 11342 3840
rect 11278 3780 11282 3836
rect 11282 3780 11338 3836
rect 11338 3780 11342 3836
rect 11278 3776 11342 3780
rect 11358 3836 11422 3840
rect 11358 3780 11362 3836
rect 11362 3780 11418 3836
rect 11418 3780 11422 3836
rect 11358 3776 11422 3780
rect 17895 3836 17959 3840
rect 17895 3780 17899 3836
rect 17899 3780 17955 3836
rect 17955 3780 17959 3836
rect 17895 3776 17959 3780
rect 17975 3836 18039 3840
rect 17975 3780 17979 3836
rect 17979 3780 18035 3836
rect 18035 3780 18039 3836
rect 17975 3776 18039 3780
rect 18055 3836 18119 3840
rect 18055 3780 18059 3836
rect 18059 3780 18115 3836
rect 18115 3780 18119 3836
rect 18055 3776 18119 3780
rect 18135 3836 18199 3840
rect 18135 3780 18139 3836
rect 18139 3780 18195 3836
rect 18195 3780 18199 3836
rect 18135 3776 18199 3780
rect 8156 3436 8220 3500
rect 7729 3292 7793 3296
rect 7729 3236 7733 3292
rect 7733 3236 7789 3292
rect 7789 3236 7793 3292
rect 7729 3232 7793 3236
rect 7809 3292 7873 3296
rect 7809 3236 7813 3292
rect 7813 3236 7869 3292
rect 7869 3236 7873 3292
rect 7809 3232 7873 3236
rect 7889 3292 7953 3296
rect 7889 3236 7893 3292
rect 7893 3236 7949 3292
rect 7949 3236 7953 3292
rect 7889 3232 7953 3236
rect 7969 3292 8033 3296
rect 7969 3236 7973 3292
rect 7973 3236 8029 3292
rect 8029 3236 8033 3292
rect 7969 3232 8033 3236
rect 14506 3292 14570 3296
rect 14506 3236 14510 3292
rect 14510 3236 14566 3292
rect 14566 3236 14570 3292
rect 14506 3232 14570 3236
rect 14586 3292 14650 3296
rect 14586 3236 14590 3292
rect 14590 3236 14646 3292
rect 14646 3236 14650 3292
rect 14586 3232 14650 3236
rect 14666 3292 14730 3296
rect 14666 3236 14670 3292
rect 14670 3236 14726 3292
rect 14726 3236 14730 3292
rect 14666 3232 14730 3236
rect 14746 3292 14810 3296
rect 14746 3236 14750 3292
rect 14750 3236 14806 3292
rect 14806 3236 14810 3292
rect 14746 3232 14810 3236
rect 4340 2748 4404 2752
rect 4340 2692 4344 2748
rect 4344 2692 4400 2748
rect 4400 2692 4404 2748
rect 4340 2688 4404 2692
rect 4420 2748 4484 2752
rect 4420 2692 4424 2748
rect 4424 2692 4480 2748
rect 4480 2692 4484 2748
rect 4420 2688 4484 2692
rect 4500 2748 4564 2752
rect 4500 2692 4504 2748
rect 4504 2692 4560 2748
rect 4560 2692 4564 2748
rect 4500 2688 4564 2692
rect 4580 2748 4644 2752
rect 4580 2692 4584 2748
rect 4584 2692 4640 2748
rect 4640 2692 4644 2748
rect 4580 2688 4644 2692
rect 11118 2748 11182 2752
rect 11118 2692 11122 2748
rect 11122 2692 11178 2748
rect 11178 2692 11182 2748
rect 11118 2688 11182 2692
rect 11198 2748 11262 2752
rect 11198 2692 11202 2748
rect 11202 2692 11258 2748
rect 11258 2692 11262 2748
rect 11198 2688 11262 2692
rect 11278 2748 11342 2752
rect 11278 2692 11282 2748
rect 11282 2692 11338 2748
rect 11338 2692 11342 2748
rect 11278 2688 11342 2692
rect 11358 2748 11422 2752
rect 11358 2692 11362 2748
rect 11362 2692 11418 2748
rect 11418 2692 11422 2748
rect 11358 2688 11422 2692
rect 17895 2748 17959 2752
rect 17895 2692 17899 2748
rect 17899 2692 17955 2748
rect 17955 2692 17959 2748
rect 17895 2688 17959 2692
rect 17975 2748 18039 2752
rect 17975 2692 17979 2748
rect 17979 2692 18035 2748
rect 18035 2692 18039 2748
rect 17975 2688 18039 2692
rect 18055 2748 18119 2752
rect 18055 2692 18059 2748
rect 18059 2692 18115 2748
rect 18115 2692 18119 2748
rect 18055 2688 18119 2692
rect 18135 2748 18199 2752
rect 18135 2692 18139 2748
rect 18139 2692 18195 2748
rect 18195 2692 18199 2748
rect 18135 2688 18199 2692
rect 7729 2204 7793 2208
rect 7729 2148 7733 2204
rect 7733 2148 7789 2204
rect 7789 2148 7793 2204
rect 7729 2144 7793 2148
rect 7809 2204 7873 2208
rect 7809 2148 7813 2204
rect 7813 2148 7869 2204
rect 7869 2148 7873 2204
rect 7809 2144 7873 2148
rect 7889 2204 7953 2208
rect 7889 2148 7893 2204
rect 7893 2148 7949 2204
rect 7949 2148 7953 2204
rect 7889 2144 7953 2148
rect 7969 2204 8033 2208
rect 7969 2148 7973 2204
rect 7973 2148 8029 2204
rect 8029 2148 8033 2204
rect 7969 2144 8033 2148
rect 14506 2204 14570 2208
rect 14506 2148 14510 2204
rect 14510 2148 14566 2204
rect 14566 2148 14570 2204
rect 14506 2144 14570 2148
rect 14586 2204 14650 2208
rect 14586 2148 14590 2204
rect 14590 2148 14646 2204
rect 14646 2148 14650 2204
rect 14586 2144 14650 2148
rect 14666 2204 14730 2208
rect 14666 2148 14670 2204
rect 14670 2148 14726 2204
rect 14726 2148 14730 2204
rect 14666 2144 14730 2148
rect 14746 2204 14810 2208
rect 14746 2148 14750 2204
rect 14750 2148 14806 2204
rect 14806 2148 14810 2204
rect 14746 2144 14810 2148
<< metal4 >>
rect 4332 22336 4653 22352
rect 4332 22272 4340 22336
rect 4404 22272 4420 22336
rect 4484 22272 4500 22336
rect 4564 22272 4580 22336
rect 4644 22272 4653 22336
rect 4332 21248 4653 22272
rect 4332 21184 4340 21248
rect 4404 21184 4420 21248
rect 4484 21184 4500 21248
rect 4564 21184 4580 21248
rect 4644 21184 4653 21248
rect 4332 20160 4653 21184
rect 4332 20096 4340 20160
rect 4404 20096 4420 20160
rect 4484 20096 4500 20160
rect 4564 20096 4580 20160
rect 4644 20096 4653 20160
rect 4332 19072 4653 20096
rect 4332 19008 4340 19072
rect 4404 19019 4420 19072
rect 4484 19019 4500 19072
rect 4564 19019 4580 19072
rect 4644 19008 4653 19072
rect 4332 18783 4374 19008
rect 4610 18783 4653 19008
rect 4332 17984 4653 18783
rect 4332 17920 4340 17984
rect 4404 17920 4420 17984
rect 4484 17920 4500 17984
rect 4564 17920 4580 17984
rect 4644 17920 4653 17984
rect 4332 16896 4653 17920
rect 4332 16832 4340 16896
rect 4404 16832 4420 16896
rect 4484 16832 4500 16896
rect 4564 16832 4580 16896
rect 4644 16832 4653 16896
rect 4332 15808 4653 16832
rect 4332 15744 4340 15808
rect 4404 15744 4420 15808
rect 4484 15744 4500 15808
rect 4564 15744 4580 15808
rect 4644 15744 4653 15808
rect 4332 14720 4653 15744
rect 4332 14656 4340 14720
rect 4404 14656 4420 14720
rect 4484 14656 4500 14720
rect 4564 14656 4580 14720
rect 4644 14656 4653 14720
rect 4332 13632 4653 14656
rect 4332 13568 4340 13632
rect 4404 13568 4420 13632
rect 4484 13568 4500 13632
rect 4564 13568 4580 13632
rect 4644 13568 4653 13632
rect 4332 12544 4653 13568
rect 4332 12480 4340 12544
rect 4404 12480 4420 12544
rect 4484 12480 4500 12544
rect 4564 12480 4580 12544
rect 4644 12480 4653 12544
rect 4332 12310 4653 12480
rect 4332 12074 4374 12310
rect 4610 12074 4653 12310
rect 4332 11456 4653 12074
rect 4332 11392 4340 11456
rect 4404 11392 4420 11456
rect 4484 11392 4500 11456
rect 4564 11392 4580 11456
rect 4644 11392 4653 11456
rect 4332 10368 4653 11392
rect 4332 10304 4340 10368
rect 4404 10304 4420 10368
rect 4484 10304 4500 10368
rect 4564 10304 4580 10368
rect 4644 10304 4653 10368
rect 4332 9280 4653 10304
rect 4332 9216 4340 9280
rect 4404 9216 4420 9280
rect 4484 9216 4500 9280
rect 4564 9216 4580 9280
rect 4644 9216 4653 9280
rect 4332 8192 4653 9216
rect 4332 8128 4340 8192
rect 4404 8128 4420 8192
rect 4484 8128 4500 8192
rect 4564 8128 4580 8192
rect 4644 8128 4653 8192
rect 4332 7104 4653 8128
rect 4332 7040 4340 7104
rect 4404 7040 4420 7104
rect 4484 7040 4500 7104
rect 4564 7040 4580 7104
rect 4644 7040 4653 7104
rect 4332 6016 4653 7040
rect 4332 5952 4340 6016
rect 4404 5952 4420 6016
rect 4484 5952 4500 6016
rect 4564 5952 4580 6016
rect 4644 5952 4653 6016
rect 4332 5600 4653 5952
rect 4332 5364 4374 5600
rect 4610 5364 4653 5600
rect 4332 4928 4653 5364
rect 4332 4864 4340 4928
rect 4404 4864 4420 4928
rect 4484 4864 4500 4928
rect 4564 4864 4580 4928
rect 4644 4864 4653 4928
rect 4332 3840 4653 4864
rect 4332 3776 4340 3840
rect 4404 3776 4420 3840
rect 4484 3776 4500 3840
rect 4564 3776 4580 3840
rect 4644 3776 4653 3840
rect 4332 2752 4653 3776
rect 4332 2688 4340 2752
rect 4404 2688 4420 2752
rect 4484 2688 4500 2752
rect 4564 2688 4580 2752
rect 4644 2688 4653 2752
rect 4332 2128 4653 2688
rect 7721 21792 8041 22352
rect 7721 21728 7729 21792
rect 7793 21728 7809 21792
rect 7873 21728 7889 21792
rect 7953 21728 7969 21792
rect 8033 21728 8041 21792
rect 7721 20704 8041 21728
rect 7721 20640 7729 20704
rect 7793 20640 7809 20704
rect 7873 20640 7889 20704
rect 7953 20640 7969 20704
rect 8033 20640 8041 20704
rect 7721 19616 8041 20640
rect 7721 19552 7729 19616
rect 7793 19552 7809 19616
rect 7873 19552 7889 19616
rect 7953 19552 7969 19616
rect 8033 19552 8041 19616
rect 7721 18528 8041 19552
rect 7721 18464 7729 18528
rect 7793 18464 7809 18528
rect 7873 18464 7889 18528
rect 7953 18464 7969 18528
rect 8033 18464 8041 18528
rect 7721 17440 8041 18464
rect 7721 17376 7729 17440
rect 7793 17376 7809 17440
rect 7873 17376 7889 17440
rect 7953 17376 7969 17440
rect 8033 17376 8041 17440
rect 7721 16352 8041 17376
rect 11110 22336 11430 22352
rect 11110 22272 11118 22336
rect 11182 22272 11198 22336
rect 11262 22272 11278 22336
rect 11342 22272 11358 22336
rect 11422 22272 11430 22336
rect 11110 21248 11430 22272
rect 11110 21184 11118 21248
rect 11182 21184 11198 21248
rect 11262 21184 11278 21248
rect 11342 21184 11358 21248
rect 11422 21184 11430 21248
rect 11110 20160 11430 21184
rect 11110 20096 11118 20160
rect 11182 20096 11198 20160
rect 11262 20096 11278 20160
rect 11342 20096 11358 20160
rect 11422 20096 11430 20160
rect 11110 19072 11430 20096
rect 11110 19008 11118 19072
rect 11182 19019 11198 19072
rect 11262 19019 11278 19072
rect 11342 19019 11358 19072
rect 11422 19008 11430 19072
rect 11110 18783 11152 19008
rect 11388 18783 11430 19008
rect 11110 17984 11430 18783
rect 11110 17920 11118 17984
rect 11182 17920 11198 17984
rect 11262 17920 11278 17984
rect 11342 17920 11358 17984
rect 11422 17920 11430 17984
rect 11110 16896 11430 17920
rect 11110 16832 11118 16896
rect 11182 16832 11198 16896
rect 11262 16832 11278 16896
rect 11342 16832 11358 16896
rect 11422 16832 11430 16896
rect 8155 16556 8221 16557
rect 8155 16492 8156 16556
rect 8220 16492 8221 16556
rect 8155 16491 8221 16492
rect 9259 16556 9325 16557
rect 9259 16492 9260 16556
rect 9324 16492 9325 16556
rect 9259 16491 9325 16492
rect 7721 16288 7729 16352
rect 7793 16288 7809 16352
rect 7873 16288 7889 16352
rect 7953 16288 7969 16352
rect 8033 16288 8041 16352
rect 7721 15664 8041 16288
rect 7721 15428 7763 15664
rect 7999 15428 8041 15664
rect 7721 15264 8041 15428
rect 7721 15200 7729 15264
rect 7793 15200 7809 15264
rect 7873 15200 7889 15264
rect 7953 15200 7969 15264
rect 8033 15200 8041 15264
rect 7721 14176 8041 15200
rect 7721 14112 7729 14176
rect 7793 14112 7809 14176
rect 7873 14112 7889 14176
rect 7953 14112 7969 14176
rect 8033 14112 8041 14176
rect 7721 13088 8041 14112
rect 7721 13024 7729 13088
rect 7793 13024 7809 13088
rect 7873 13024 7889 13088
rect 7953 13024 7969 13088
rect 8033 13024 8041 13088
rect 7721 12000 8041 13024
rect 8158 12477 8218 16491
rect 9262 14109 9322 16491
rect 11110 15808 11430 16832
rect 11110 15744 11118 15808
rect 11182 15744 11198 15808
rect 11262 15744 11278 15808
rect 11342 15744 11358 15808
rect 11422 15744 11430 15808
rect 11110 14720 11430 15744
rect 11110 14656 11118 14720
rect 11182 14656 11198 14720
rect 11262 14656 11278 14720
rect 11342 14656 11358 14720
rect 11422 14656 11430 14720
rect 9259 14108 9325 14109
rect 9259 14044 9260 14108
rect 9324 14044 9325 14108
rect 9259 14043 9325 14044
rect 11110 13632 11430 14656
rect 11110 13568 11118 13632
rect 11182 13568 11198 13632
rect 11262 13568 11278 13632
rect 11342 13568 11358 13632
rect 11422 13568 11430 13632
rect 11110 12544 11430 13568
rect 11110 12480 11118 12544
rect 11182 12480 11198 12544
rect 11262 12480 11278 12544
rect 11342 12480 11358 12544
rect 11422 12480 11430 12544
rect 8155 12476 8221 12477
rect 8155 12412 8156 12476
rect 8220 12412 8221 12476
rect 8155 12411 8221 12412
rect 7721 11936 7729 12000
rect 7793 11936 7809 12000
rect 7873 11936 7889 12000
rect 7953 11936 7969 12000
rect 8033 11936 8041 12000
rect 7721 10912 8041 11936
rect 7721 10848 7729 10912
rect 7793 10848 7809 10912
rect 7873 10848 7889 10912
rect 7953 10848 7969 10912
rect 8033 10848 8041 10912
rect 7721 9824 8041 10848
rect 7721 9760 7729 9824
rect 7793 9760 7809 9824
rect 7873 9760 7889 9824
rect 7953 9760 7969 9824
rect 8033 9760 8041 9824
rect 7721 8955 8041 9760
rect 7721 8736 7763 8955
rect 7999 8736 8041 8955
rect 7721 8672 7729 8736
rect 7793 8672 7809 8719
rect 7873 8672 7889 8719
rect 7953 8672 7969 8719
rect 8033 8672 8041 8736
rect 7721 7648 8041 8672
rect 7721 7584 7729 7648
rect 7793 7584 7809 7648
rect 7873 7584 7889 7648
rect 7953 7584 7969 7648
rect 8033 7584 8041 7648
rect 7721 6560 8041 7584
rect 11110 12310 11430 12480
rect 11110 12074 11152 12310
rect 11388 12074 11430 12310
rect 11110 11456 11430 12074
rect 11110 11392 11118 11456
rect 11182 11392 11198 11456
rect 11262 11392 11278 11456
rect 11342 11392 11358 11456
rect 11422 11392 11430 11456
rect 11110 10368 11430 11392
rect 11110 10304 11118 10368
rect 11182 10304 11198 10368
rect 11262 10304 11278 10368
rect 11342 10304 11358 10368
rect 11422 10304 11430 10368
rect 11110 9280 11430 10304
rect 11110 9216 11118 9280
rect 11182 9216 11198 9280
rect 11262 9216 11278 9280
rect 11342 9216 11358 9280
rect 11422 9216 11430 9280
rect 11110 8192 11430 9216
rect 11110 8128 11118 8192
rect 11182 8128 11198 8192
rect 11262 8128 11278 8192
rect 11342 8128 11358 8192
rect 11422 8128 11430 8192
rect 11110 7104 11430 8128
rect 11110 7040 11118 7104
rect 11182 7040 11198 7104
rect 11262 7040 11278 7104
rect 11342 7040 11358 7104
rect 11422 7040 11430 7104
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 7721 6496 7729 6560
rect 7793 6496 7809 6560
rect 7873 6496 7889 6560
rect 7953 6496 7969 6560
rect 8033 6496 8041 6560
rect 7721 5472 8041 6496
rect 7721 5408 7729 5472
rect 7793 5408 7809 5472
rect 7873 5408 7889 5472
rect 7953 5408 7969 5472
rect 8033 5408 8041 5472
rect 7721 4384 8041 5408
rect 7721 4320 7729 4384
rect 7793 4320 7809 4384
rect 7873 4320 7889 4384
rect 7953 4320 7969 4384
rect 8033 4320 8041 4384
rect 7721 3296 8041 4320
rect 8158 3501 8218 6971
rect 11110 6016 11430 7040
rect 11110 5952 11118 6016
rect 11182 5952 11198 6016
rect 11262 5952 11278 6016
rect 11342 5952 11358 6016
rect 11422 5952 11430 6016
rect 11110 5600 11430 5952
rect 9443 5404 9509 5405
rect 9443 5340 9444 5404
rect 9508 5340 9509 5404
rect 9443 5339 9509 5340
rect 11110 5364 11152 5600
rect 11388 5364 11430 5600
rect 9446 4861 9506 5339
rect 11110 4928 11430 5364
rect 11110 4864 11118 4928
rect 11182 4864 11198 4928
rect 11262 4864 11278 4928
rect 11342 4864 11358 4928
rect 11422 4864 11430 4928
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 11110 3840 11430 4864
rect 11110 3776 11118 3840
rect 11182 3776 11198 3840
rect 11262 3776 11278 3840
rect 11342 3776 11358 3840
rect 11422 3776 11430 3840
rect 8155 3500 8221 3501
rect 8155 3436 8156 3500
rect 8220 3436 8221 3500
rect 8155 3435 8221 3436
rect 7721 3232 7729 3296
rect 7793 3232 7809 3296
rect 7873 3232 7889 3296
rect 7953 3232 7969 3296
rect 8033 3232 8041 3296
rect 7721 2208 8041 3232
rect 7721 2144 7729 2208
rect 7793 2144 7809 2208
rect 7873 2144 7889 2208
rect 7953 2144 7969 2208
rect 8033 2144 8041 2208
rect 7721 2128 8041 2144
rect 11110 2752 11430 3776
rect 11110 2688 11118 2752
rect 11182 2688 11198 2752
rect 11262 2688 11278 2752
rect 11342 2688 11358 2752
rect 11422 2688 11430 2752
rect 11110 2128 11430 2688
rect 14498 21792 14818 22352
rect 14498 21728 14506 21792
rect 14570 21728 14586 21792
rect 14650 21728 14666 21792
rect 14730 21728 14746 21792
rect 14810 21728 14818 21792
rect 14498 20704 14818 21728
rect 14498 20640 14506 20704
rect 14570 20640 14586 20704
rect 14650 20640 14666 20704
rect 14730 20640 14746 20704
rect 14810 20640 14818 20704
rect 14498 19616 14818 20640
rect 14498 19552 14506 19616
rect 14570 19552 14586 19616
rect 14650 19552 14666 19616
rect 14730 19552 14746 19616
rect 14810 19552 14818 19616
rect 14498 18528 14818 19552
rect 17887 22336 18207 22352
rect 17887 22272 17895 22336
rect 17959 22272 17975 22336
rect 18039 22272 18055 22336
rect 18119 22272 18135 22336
rect 18199 22272 18207 22336
rect 17887 21248 18207 22272
rect 17887 21184 17895 21248
rect 17959 21184 17975 21248
rect 18039 21184 18055 21248
rect 18119 21184 18135 21248
rect 18199 21184 18207 21248
rect 17887 20160 18207 21184
rect 20299 20772 20365 20773
rect 20299 20708 20300 20772
rect 20364 20708 20365 20772
rect 20299 20707 20365 20708
rect 20483 20772 20549 20773
rect 20483 20708 20484 20772
rect 20548 20708 20549 20772
rect 20483 20707 20549 20708
rect 17887 20096 17895 20160
rect 17959 20096 17975 20160
rect 18039 20096 18055 20160
rect 18119 20096 18135 20160
rect 18199 20096 18207 20160
rect 14963 19276 15029 19277
rect 14963 19212 14964 19276
rect 15028 19212 15029 19276
rect 14963 19211 15029 19212
rect 14498 18464 14506 18528
rect 14570 18464 14586 18528
rect 14650 18464 14666 18528
rect 14730 18464 14746 18528
rect 14810 18464 14818 18528
rect 14498 17440 14818 18464
rect 14498 17376 14506 17440
rect 14570 17376 14586 17440
rect 14650 17376 14666 17440
rect 14730 17376 14746 17440
rect 14810 17376 14818 17440
rect 14498 16352 14818 17376
rect 14498 16288 14506 16352
rect 14570 16288 14586 16352
rect 14650 16288 14666 16352
rect 14730 16288 14746 16352
rect 14810 16288 14818 16352
rect 14498 15664 14818 16288
rect 14498 15428 14540 15664
rect 14776 15428 14818 15664
rect 14498 15264 14818 15428
rect 14498 15200 14506 15264
rect 14570 15200 14586 15264
rect 14650 15200 14666 15264
rect 14730 15200 14746 15264
rect 14810 15200 14818 15264
rect 14498 14176 14818 15200
rect 14498 14112 14506 14176
rect 14570 14112 14586 14176
rect 14650 14112 14666 14176
rect 14730 14112 14746 14176
rect 14810 14112 14818 14176
rect 14498 13088 14818 14112
rect 14966 13429 15026 19211
rect 17887 19072 18207 20096
rect 19931 19684 19997 19685
rect 19931 19620 19932 19684
rect 19996 19620 19997 19684
rect 19931 19619 19997 19620
rect 17887 19008 17895 19072
rect 17959 19019 17975 19072
rect 18039 19019 18055 19072
rect 18119 19019 18135 19072
rect 18199 19008 18207 19072
rect 17887 18783 17929 19008
rect 18165 18783 18207 19008
rect 17887 17984 18207 18783
rect 17887 17920 17895 17984
rect 17959 17920 17975 17984
rect 18039 17920 18055 17984
rect 18119 17920 18135 17984
rect 18199 17920 18207 17984
rect 17887 16896 18207 17920
rect 17887 16832 17895 16896
rect 17959 16832 17975 16896
rect 18039 16832 18055 16896
rect 18119 16832 18135 16896
rect 18199 16832 18207 16896
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17726 13973 17786 16627
rect 17887 15808 18207 16832
rect 17887 15744 17895 15808
rect 17959 15744 17975 15808
rect 18039 15744 18055 15808
rect 18119 15744 18135 15808
rect 18199 15744 18207 15808
rect 17887 14720 18207 15744
rect 17887 14656 17895 14720
rect 17959 14656 17975 14720
rect 18039 14656 18055 14720
rect 18119 14656 18135 14720
rect 18199 14656 18207 14720
rect 17723 13972 17789 13973
rect 17723 13908 17724 13972
rect 17788 13908 17789 13972
rect 17723 13907 17789 13908
rect 17887 13632 18207 14656
rect 17887 13568 17895 13632
rect 17959 13568 17975 13632
rect 18039 13568 18055 13632
rect 18119 13568 18135 13632
rect 18199 13568 18207 13632
rect 14963 13428 15029 13429
rect 14963 13364 14964 13428
rect 15028 13364 15029 13428
rect 14963 13363 15029 13364
rect 14498 13024 14506 13088
rect 14570 13024 14586 13088
rect 14650 13024 14666 13088
rect 14730 13024 14746 13088
rect 14810 13024 14818 13088
rect 14498 12000 14818 13024
rect 14498 11936 14506 12000
rect 14570 11936 14586 12000
rect 14650 11936 14666 12000
rect 14730 11936 14746 12000
rect 14810 11936 14818 12000
rect 14498 10912 14818 11936
rect 14498 10848 14506 10912
rect 14570 10848 14586 10912
rect 14650 10848 14666 10912
rect 14730 10848 14746 10912
rect 14810 10848 14818 10912
rect 14498 9824 14818 10848
rect 14498 9760 14506 9824
rect 14570 9760 14586 9824
rect 14650 9760 14666 9824
rect 14730 9760 14746 9824
rect 14810 9760 14818 9824
rect 14498 8955 14818 9760
rect 14498 8736 14540 8955
rect 14776 8736 14818 8955
rect 14498 8672 14506 8736
rect 14570 8672 14586 8719
rect 14650 8672 14666 8719
rect 14730 8672 14746 8719
rect 14810 8672 14818 8736
rect 14498 7648 14818 8672
rect 14498 7584 14506 7648
rect 14570 7584 14586 7648
rect 14650 7584 14666 7648
rect 14730 7584 14746 7648
rect 14810 7584 14818 7648
rect 14498 6560 14818 7584
rect 14498 6496 14506 6560
rect 14570 6496 14586 6560
rect 14650 6496 14666 6560
rect 14730 6496 14746 6560
rect 14810 6496 14818 6560
rect 14498 5472 14818 6496
rect 14498 5408 14506 5472
rect 14570 5408 14586 5472
rect 14650 5408 14666 5472
rect 14730 5408 14746 5472
rect 14810 5408 14818 5472
rect 14498 4384 14818 5408
rect 14498 4320 14506 4384
rect 14570 4320 14586 4384
rect 14650 4320 14666 4384
rect 14730 4320 14746 4384
rect 14810 4320 14818 4384
rect 14498 3296 14818 4320
rect 14498 3232 14506 3296
rect 14570 3232 14586 3296
rect 14650 3232 14666 3296
rect 14730 3232 14746 3296
rect 14810 3232 14818 3296
rect 14498 2208 14818 3232
rect 14498 2144 14506 2208
rect 14570 2144 14586 2208
rect 14650 2144 14666 2208
rect 14730 2144 14746 2208
rect 14810 2144 14818 2208
rect 14498 2128 14818 2144
rect 17887 12544 18207 13568
rect 17887 12480 17895 12544
rect 17959 12480 17975 12544
rect 18039 12480 18055 12544
rect 18119 12480 18135 12544
rect 18199 12480 18207 12544
rect 17887 12310 18207 12480
rect 17887 12074 17929 12310
rect 18165 12074 18207 12310
rect 17887 11456 18207 12074
rect 17887 11392 17895 11456
rect 17959 11392 17975 11456
rect 18039 11392 18055 11456
rect 18119 11392 18135 11456
rect 18199 11392 18207 11456
rect 17887 10368 18207 11392
rect 17887 10304 17895 10368
rect 17959 10304 17975 10368
rect 18039 10304 18055 10368
rect 18119 10304 18135 10368
rect 18199 10304 18207 10368
rect 17887 9280 18207 10304
rect 17887 9216 17895 9280
rect 17959 9216 17975 9280
rect 18039 9216 18055 9280
rect 18119 9216 18135 9280
rect 18199 9216 18207 9280
rect 17887 8192 18207 9216
rect 19934 9077 19994 19619
rect 20115 19548 20181 19549
rect 20115 19484 20116 19548
rect 20180 19484 20181 19548
rect 20115 19483 20181 19484
rect 19931 9076 19997 9077
rect 19931 9012 19932 9076
rect 19996 9012 19997 9076
rect 19931 9011 19997 9012
rect 17887 8128 17895 8192
rect 17959 8128 17975 8192
rect 18039 8128 18055 8192
rect 18119 8128 18135 8192
rect 18199 8128 18207 8192
rect 17887 7104 18207 8128
rect 17887 7040 17895 7104
rect 17959 7040 17975 7104
rect 18039 7040 18055 7104
rect 18119 7040 18135 7104
rect 18199 7040 18207 7104
rect 17887 6016 18207 7040
rect 17887 5952 17895 6016
rect 17959 5952 17975 6016
rect 18039 5952 18055 6016
rect 18119 5952 18135 6016
rect 18199 5952 18207 6016
rect 17887 5600 18207 5952
rect 20118 5949 20178 19483
rect 20302 9485 20362 20707
rect 20299 9484 20365 9485
rect 20299 9420 20300 9484
rect 20364 9420 20365 9484
rect 20299 9419 20365 9420
rect 20486 7445 20546 20707
rect 20483 7444 20549 7445
rect 20483 7380 20484 7444
rect 20548 7380 20549 7444
rect 20483 7379 20549 7380
rect 20115 5948 20181 5949
rect 20115 5884 20116 5948
rect 20180 5884 20181 5948
rect 20115 5883 20181 5884
rect 17887 5364 17929 5600
rect 18165 5364 18207 5600
rect 17887 4928 18207 5364
rect 17887 4864 17895 4928
rect 17959 4864 17975 4928
rect 18039 4864 18055 4928
rect 18119 4864 18135 4928
rect 18199 4864 18207 4928
rect 17887 3840 18207 4864
rect 17887 3776 17895 3840
rect 17959 3776 17975 3840
rect 18039 3776 18055 3840
rect 18119 3776 18135 3840
rect 18199 3776 18207 3840
rect 17887 2752 18207 3776
rect 17887 2688 17895 2752
rect 17959 2688 17975 2752
rect 18039 2688 18055 2752
rect 18119 2688 18135 2752
rect 18199 2688 18207 2752
rect 17887 2128 18207 2688
<< via4 >>
rect 4374 19008 4404 19019
rect 4404 19008 4420 19019
rect 4420 19008 4484 19019
rect 4484 19008 4500 19019
rect 4500 19008 4564 19019
rect 4564 19008 4580 19019
rect 4580 19008 4610 19019
rect 4374 18783 4610 19008
rect 4374 12074 4610 12310
rect 4374 5364 4610 5600
rect 11152 19008 11182 19019
rect 11182 19008 11198 19019
rect 11198 19008 11262 19019
rect 11262 19008 11278 19019
rect 11278 19008 11342 19019
rect 11342 19008 11358 19019
rect 11358 19008 11388 19019
rect 11152 18783 11388 19008
rect 7763 15428 7999 15664
rect 7763 8736 7999 8955
rect 7763 8719 7793 8736
rect 7793 8719 7809 8736
rect 7809 8719 7873 8736
rect 7873 8719 7889 8736
rect 7889 8719 7953 8736
rect 7953 8719 7969 8736
rect 7969 8719 7999 8736
rect 11152 12074 11388 12310
rect 11152 5364 11388 5600
rect 14540 15428 14776 15664
rect 17929 19008 17959 19019
rect 17959 19008 17975 19019
rect 17975 19008 18039 19019
rect 18039 19008 18055 19019
rect 18055 19008 18119 19019
rect 18119 19008 18135 19019
rect 18135 19008 18165 19019
rect 17929 18783 18165 19008
rect 14540 8736 14776 8955
rect 14540 8719 14570 8736
rect 14570 8719 14586 8736
rect 14586 8719 14650 8736
rect 14650 8719 14666 8736
rect 14666 8719 14730 8736
rect 14730 8719 14746 8736
rect 14746 8719 14776 8736
rect 17929 12074 18165 12310
rect 17929 5364 18165 5600
<< metal5 >>
rect 1104 19019 21436 19061
rect 1104 18783 4374 19019
rect 4610 18783 11152 19019
rect 11388 18783 17929 19019
rect 18165 18783 21436 19019
rect 1104 18741 21436 18783
rect 1104 15664 21436 15706
rect 1104 15428 7763 15664
rect 7999 15428 14540 15664
rect 14776 15428 21436 15664
rect 1104 15386 21436 15428
rect 1104 12310 21436 12352
rect 1104 12074 4374 12310
rect 4610 12074 11152 12310
rect 11388 12074 17929 12310
rect 18165 12074 21436 12310
rect 1104 12032 21436 12074
rect 1104 8955 21436 8997
rect 1104 8719 7763 8955
rect 7999 8719 14540 8955
rect 14776 8719 21436 8955
rect 1104 8677 21436 8719
rect 1104 5600 21436 5643
rect 1104 5364 4374 5600
rect 4610 5364 11152 5600
rect 11388 5364 17929 5600
rect 18165 5364 21436 5600
rect 1104 5322 21436 5364
use sky130_fd_sc_hd__clkbuf_2  input15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0949_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 1472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1632469394
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1632469394
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1632469394
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1632469394
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1632469394
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1632469394
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1632469394
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 1632469394
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1632469394
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1632469394
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37
timestamp 1632469394
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1632469394
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp 1632469394
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 5060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _0820_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3680 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1632469394
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0812_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 5244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1632469394
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1632469394
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1632469394
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1632469394
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 6624 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1632469394
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1632469394
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1632469394
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1632469394
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1632469394
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1632469394
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1632469394
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73
timestamp 1632469394
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1632469394
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1632469394
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1632469394
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1632469394
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1632469394
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9016 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1632469394
transform 1 0 7820 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1632469394
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1632469394
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1632469394
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97
timestamp 1632469394
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1632469394
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1632469394
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_97
timestamp 1632469394
transform 1 0 10028 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 10120 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1632469394
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 10120 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1632469394
transform 1 0 11868 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 12052 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1632469394
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1632469394
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1632469394
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1632469394
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1632469394
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1632469394
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1632469394
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1632469394
transform 1 0 13156 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1632469394
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1632469394
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1632469394
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1632469394
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_140
timestamp 1632469394
transform 1 0 13984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1632469394
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1632469394
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1632469394
transform 1 0 14076 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1632469394
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1632469394
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1632469394
transform 1 0 15272 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1632469394
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1632469394
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1632469394
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1632469394
transform 1 0 16652 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 16744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1632469394
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1632469394
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1632469394
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1632469394
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1632469394
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1632469394
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1632469394
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1632469394
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1632469394
transform 1 0 17296 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1632469394
transform 1 0 17848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_191
timestamp 1632469394
transform 1 0 18676 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1632469394
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1632469394
transform 1 0 17940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1632469394
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1632469394
transform 1 0 19228 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_1_205
timestamp 1632469394
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1632469394
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1632469394
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1632469394
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 20516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1632469394
transform -1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1632469394
transform -1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_217
timestamp 1632469394
transform 1 0 21068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1632469394
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1632469394
transform 1 0 20792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_11
timestamp 1632469394
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1632469394
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1632469394
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1632469394
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1632469394
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1632469394
transform 1 0 2944 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1632469394
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1632469394
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1632469394
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1632469394
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0818_
timestamp 1632469394
transform 1 0 3864 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1632469394
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1632469394
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1632469394
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 6716 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1632469394
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1632469394
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1632469394
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1632469394
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0815_
timestamp 1632469394
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1632469394
transform 1 0 11132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1632469394
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0914_
timestamp 1632469394
transform 1 0 9292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0932_
timestamp 1632469394
transform 1 0 10396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1632469394
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_127
timestamp 1632469394
transform 1 0 12788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _0896_
timestamp 1632469394
transform 1 0 12880 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0904_
timestamp 1632469394
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1632469394
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1632469394
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1632469394
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _0897_
timestamp 1632469394
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1632469394
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_164
timestamp 1632469394
transform 1 0 16192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_169
timestamp 1632469394
transform 1 0 16652 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0862_
timestamp 1632469394
transform 1 0 15180 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 1632469394
transform 1 0 17020 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1632469394
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1632469394
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1632469394
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1632469394
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 19504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1632469394
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_206
timestamp 1632469394
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1632469394
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1632469394
transform -1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1632469394
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1632469394
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1632469394
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1632469394
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1632469394
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1632469394
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1632469394
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1632469394
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1632469394
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1632469394
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1632469394
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3864 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1632469394
transform 1 0 4876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1632469394
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1632469394
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1632469394
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1632469394
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1632469394
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1632469394
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1632469394
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1632469394
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0918_
timestamp 1632469394
transform 1 0 8372 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1632469394
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1632469394
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1632469394
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1632469394
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0925_
timestamp 1632469394
transform 1 0 9476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1632469394
transform 1 0 10672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1632469394
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1632469394
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1632469394
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0905_
timestamp 1632469394
transform 1 0 12604 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _0906_
timestamp 1632469394
transform 1 0 11592 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1632469394
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_140
timestamp 1632469394
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1632469394
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1632469394
transform 1 0 14536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1632469394
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1632469394
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1632469394
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_174
timestamp 1632469394
transform 1 0 17112 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1632469394
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 16652 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0861_
timestamp 1632469394
transform 1 0 15272 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1632469394
transform 1 0 17848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1632469394
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1632469394
transform 1 0 17940 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1632469394
transform 1 0 18768 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1632469394
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1632469394
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1632469394
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_214
timestamp 1632469394
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1632469394
transform -1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1632469394
transform 1 0 19780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1632469394
transform 1 0 20424 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1632469394
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1632469394
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1632469394
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1632469394
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1632469394
transform 1 0 1380 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1632469394
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1632469394
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1632469394
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0831_
timestamp 1632469394
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1632469394
transform 1 0 5152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1632469394
transform 1 0 5888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59
timestamp 1632469394
transform 1 0 6532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0826_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 5980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1632469394
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_69
timestamp 1632469394
transform 1 0 7452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_75
timestamp 1632469394
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1632469394
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1632469394
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _0927_
timestamp 1632469394
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1632469394
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1632469394
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_92
timestamp 1632469394
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1632469394
transform 1 0 10948 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9936 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1632469394
transform 1 0 11408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1632469394
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1632469394
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0917_
timestamp 1632469394
transform 1 0 11776 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1632469394
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1632469394
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1632469394
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1632469394
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1632469394
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1632469394
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1632469394
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_167
timestamp 1632469394
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0835_
timestamp 1632469394
transform 1 0 15916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0853_
timestamp 1632469394
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1632469394
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1632469394
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1632469394
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1632469394
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1632469394
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1632469394
transform 1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0859_
timestamp 1632469394
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1632469394
transform 1 0 19964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1632469394
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1632469394
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1632469394
transform -1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1632469394
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_11
timestamp 1632469394
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1632469394
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1632469394
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_4  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 2852 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1632469394
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1632469394
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _0829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 4784 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1632469394
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1632469394
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_61
timestamp 1632469394
transform 1 0 6716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1632469394
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0827_
timestamp 1632469394
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_74
timestamp 1632469394
transform 1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1632469394
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1632469394
transform 1 0 9108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0833_
timestamp 1632469394
transform 1 0 7268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1632469394
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1632469394
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1632469394
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1632469394
transform 1 0 10672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp 1632469394
transform 1 0 9476 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1632469394
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 1632469394
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_126
timestamp 1632469394
transform 1 0 12696 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1632469394
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0903_
timestamp 1632469394
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0944_
timestamp 1632469394
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1632469394
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_152
timestamp 1632469394
transform 1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _0899_
timestamp 1632469394
transform 1 0 14444 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1632469394
transform 1 0 13248 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1632469394
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1632469394
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1632469394
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1632469394
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1632469394
transform 1 0 17480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1632469394
transform 1 0 17848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1632469394
transform 1 0 18308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 18676 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1632469394
transform 1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_198
timestamp 1632469394
transform 1 0 19320 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1632469394
transform 1 0 19872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_212
timestamp 1632469394
transform 1 0 20608 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1632469394
transform -1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0848_
timestamp 1632469394
transform 1 0 19964 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1632469394
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1632469394
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1632469394
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1632469394
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1632469394
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1632469394
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0808_
timestamp 1632469394
transform 1 0 2024 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_6_11
timestamp 1632469394
transform 1 0 2116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0841_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1632469394
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1632469394
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1632469394
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_43
timestamp 1632469394
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1632469394
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_37
timestamp 1632469394
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1632469394
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0843_
timestamp 1632469394
transform 1 0 4324 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0844_
timestamp 1632469394
transform 1 0 4876 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_51
timestamp 1632469394
transform 1 0 5796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_61
timestamp 1632469394
transform 1 0 6716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1632469394
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1632469394
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1632469394
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_64
timestamp 1632469394
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1632469394
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0828_
timestamp 1632469394
transform 1 0 6440 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1632469394
transform 1 0 5888 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1632469394
transform 1 0 7360 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1632469394
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_71
timestamp 1632469394
transform 1 0 7636 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1632469394
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0958_
timestamp 1632469394
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1632469394
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1632469394
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1632469394
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1632469394
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1632469394
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1632469394
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1632469394
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 1632469394
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1632469394
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1632469394
transform 1 0 10304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_104
timestamp 1632469394
transform 1 0 10672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1632469394
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1632469394
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0923_
timestamp 1632469394
transform 1 0 9200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1632469394
transform 1 0 9476 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp 1632469394
transform 1 0 10120 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1632469394
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1632469394
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_119
timestamp 1632469394
transform 1 0 12052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_128
timestamp 1632469394
transform 1 0 12880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1632469394
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1632469394
transform 1 0 12420 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1632469394
transform 1 0 11316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0913_
timestamp 1632469394
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1632469394
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1632469394
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_147
timestamp 1632469394
transform 1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1632469394
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1632469394
transform 1 0 14628 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1632469394
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0886_
timestamp 1632469394
transform 1 0 14168 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1632469394
transform 1 0 13248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0890_
timestamp 1632469394
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1632469394
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0850_
timestamp 1632469394
transform 1 0 15548 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1632469394
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_157
timestamp 1632469394
transform 1 0 15548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1632469394
transform 1 0 16100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1632469394
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1632469394
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1632469394
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_169
timestamp 1632469394
transform 1 0 16652 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_172
timestamp 1632469394
transform 1 0 16928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1632469394
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1632469394
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1632469394
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_180
timestamp 1632469394
transform 1 0 17664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1632469394
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 18216 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_4  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 17756 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1632469394
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1632469394
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_214
timestamp 1632469394
transform 1 0 20792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_202
timestamp 1632469394
transform 1 0 19688 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_214
timestamp 1632469394
transform 1 0 20792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1632469394
transform -1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1632469394
transform -1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 1632469394
transform 1 0 19964 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1632469394
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1632469394
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1632469394
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1632469394
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1632469394
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1632469394
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1632469394
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 1632469394
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1632469394
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_33
timestamp 1632469394
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1632469394
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1632469394
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1632469394
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_47
timestamp 1632469394
transform 1 0 5428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1632469394
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0810_
timestamp 1632469394
transform 1 0 5980 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1632469394
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1632469394
transform 1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_67
timestamp 1632469394
transform 1 0 7268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1632469394
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1632469394
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_1  _0832_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 7820 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1632469394
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1632469394
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1632469394
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1632469394
transform 1 0 9568 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0924_
timestamp 1632469394
transform 1 0 10580 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1632469394
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1632469394
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1632469394
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0902_
timestamp 1632469394
transform 1 0 12512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1632469394
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1632469394
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1632469394
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1632469394
transform 1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1632469394
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_1  _0849_
timestamp 1632469394
transform 1 0 14812 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1632469394
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1632469394
transform 1 0 14168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1632469394
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_166
timestamp 1632469394
transform 1 0 16376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1632469394
transform 1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0501_
timestamp 1632469394
transform 1 0 15824 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1632469394
transform 1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp 1632469394
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1632469394
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1632469394
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1632469394
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1632469394
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0882_
timestamp 1632469394
transform 1 0 18124 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1632469394
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_211
timestamp 1632469394
transform 1 0 20516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_217
timestamp 1632469394
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1632469394
transform -1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0872_
timestamp 1632469394
transform 1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_11
timestamp 1632469394
transform 1 0 2116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1632469394
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1632469394
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1632469394
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1632469394
transform 1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1632469394
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1632469394
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_37
timestamp 1632469394
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_2  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3588 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_9_45
timestamp 1632469394
transform 1 0 5244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1632469394
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1632469394
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1632469394
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0809_
timestamp 1632469394
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_66
timestamp 1632469394
transform 1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_74
timestamp 1632469394
transform 1 0 7912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1632469394
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0498_
timestamp 1632469394
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1632469394
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_100
timestamp 1632469394
transform 1 0 10304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_104
timestamp 1632469394
transform 1 0 10672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1632469394
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1632469394
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1632469394
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_1  _0919_
timestamp 1632469394
transform 1 0 9660 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1632469394
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_119
timestamp 1632469394
transform 1 0 12052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1632469394
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_130
timestamp 1632469394
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1632469394
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0500_
timestamp 1632469394
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0822_
timestamp 1632469394
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_141
timestamp 1632469394
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_147
timestamp 1632469394
transform 1 0 14628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1632469394
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _0898_
timestamp 1632469394
transform 1 0 13432 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1632469394
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1632469394
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1632469394
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0873_
timestamp 1632469394
transform 1 0 15364 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_1  _0874_
timestamp 1632469394
transform 1 0 16652 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_176
timestamp 1632469394
transform 1 0 17296 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_191
timestamp 1632469394
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1632469394
transform 1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1632469394
transform 1 0 19044 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1632469394
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_204
timestamp 1632469394
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1632469394
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1632469394
transform -1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1632469394
transform 1 0 19964 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1632469394
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1632469394
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1632469394
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1632469394
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0805_
timestamp 1632469394
transform 1 0 2300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1632469394
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1632469394
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_39
timestamp 1632469394
transform 1 0 4692 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1632469394
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1632469394
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1632469394
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1632469394
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_50
timestamp 1632469394
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_57
timestamp 1632469394
transform 1 0 6348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1632469394
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _0798_
timestamp 1632469394
transform 1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1632469394
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1632469394
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1632469394
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1632469394
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp 1632469394
transform 1 0 7268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_104
timestamp 1632469394
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1632469394
transform 1 0 9200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0920_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1632469394
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_111
timestamp 1632469394
transform 1 0 11316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1632469394
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _0907_
timestamp 1632469394
transform 1 0 11868 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0908_
timestamp 1632469394
transform 1 0 12880 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1632469394
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1632469394
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1632469394
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1632469394
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1632469394
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1632469394
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0497_
timestamp 1632469394
transform 1 0 14536 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_161
timestamp 1632469394
transform 1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_169
timestamp 1632469394
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1632469394
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1632469394
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _0885_
timestamp 1632469394
transform 1 0 15272 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1632469394
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1632469394
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1632469394
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1632469394
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 18124 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_205
timestamp 1632469394
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1632469394
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_214
timestamp 1632469394
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1632469394
transform -1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0883_
timestamp 1632469394
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1632469394
transform 1 0 20424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1632469394
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1632469394
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1632469394
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1632469394
transform 1 0 2668 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _0792_
timestamp 1632469394
transform 1 0 1656 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1632469394
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_36
timestamp 1632469394
transform 1 0 4416 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1007_
timestamp 1632469394
transform 1 0 4968 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1632469394
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1632469394
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1632469394
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1632469394
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0794_
timestamp 1632469394
transform 1 0 6716 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_70
timestamp 1632469394
transform 1 0 7544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1632469394
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _0935_
timestamp 1632469394
transform 1 0 8280 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1632469394
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1632469394
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1632469394
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0502_
timestamp 1632469394
transform 1 0 10488 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1632469394
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1632469394
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1632469394
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1632469394
transform 1 0 12052 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1632469394
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_144
timestamp 1632469394
transform 1 0 14352 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0512_
timestamp 1632469394
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0799_
timestamp 1632469394
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1632469394
transform 1 0 15088 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1632469394
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1632469394
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1632469394
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1632469394
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0878_
timestamp 1632469394
transform 1 0 16928 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1632469394
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1632469394
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1632469394
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1632469394
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0870_
timestamp 1632469394
transform 1 0 19136 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1632469394
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_203
timestamp 1632469394
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_210
timestamp 1632469394
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1632469394
transform -1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1632469394
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_11
timestamp 1632469394
transform 1 0 2116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1632469394
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1632469394
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1632469394
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1632469394
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1632469394
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1632469394
transform 1 0 4048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1632469394
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1632469394
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1632469394
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp 1632469394
transform 1 0 4508 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1632469394
transform 1 0 5336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1632469394
transform 1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _0795_
timestamp 1632469394
transform 1 0 6992 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0800_
timestamp 1632469394
transform 1 0 5704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_71
timestamp 1632469394
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1632469394
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1632469394
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1632469394
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1632469394
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0793_
timestamp 1632469394
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_88
timestamp 1632469394
transform 1 0 9200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_94
timestamp 1632469394
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_4  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9844 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1632469394
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1632469394
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_128
timestamp 1632469394
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0510_
timestamp 1632469394
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0776_
timestamp 1632469394
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1632469394
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1632469394
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1632469394
transform 1 0 14444 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1632469394
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0814_
timestamp 1632469394
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_162
timestamp 1632469394
transform 1 0 16008 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1632469394
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0867_
timestamp 1632469394
transform 1 0 16652 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0884_
timestamp 1632469394
transform 1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_175
timestamp 1632469394
transform 1 0 17204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_188
timestamp 1632469394
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1632469394
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1632469394
transform 1 0 17572 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_206
timestamp 1632469394
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_214
timestamp 1632469394
transform 1 0 20792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1632469394
transform -1 0 21436 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1632469394
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1632469394
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1632469394
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1632469394
transform 1 0 1472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1632469394
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1632469394
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1632469394
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1632469394
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1632469394
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0791_
timestamp 1632469394
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0775_
timestamp 1632469394
transform 1 0 2300 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1632469394
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1632469394
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1632469394
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1632469394
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1632469394
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1632469394
transform 1 0 3864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1632469394
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1632469394
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1632469394
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1632469394
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0780_
timestamp 1632469394
transform 1 0 4692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_33
timestamp 1632469394
transform 1 0 4140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_31
timestamp 1632469394
transform 1 0 3956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_40
timestamp 1632469394
transform 1 0 4784 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1632469394
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1632469394
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_60
timestamp 1632469394
transform 1 0 6624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_49
timestamp 1632469394
transform 1 0 5612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_57
timestamp 1632469394
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1632469394
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 1632469394
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1632469394
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0797_
timestamp 1632469394
transform 1 0 5428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1632469394
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0782_
timestamp 1632469394
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1632469394
transform 1 0 8004 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1632469394
transform 1 0 7268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1632469394
transform 1 0 7820 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1632469394
transform 1 0 7360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1632469394
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1632469394
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1632469394
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1632469394
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1632469394
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_8  _0999_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 8648 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1632469394
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1632469394
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_94
timestamp 1632469394
transform 1 0 9752 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0929_
timestamp 1632469394
transform 1 0 10304 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0685_
timestamp 1632469394
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0523_
timestamp 1632469394
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1632469394
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1632469394
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0662_
timestamp 1632469394
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1632469394
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_117
timestamp 1632469394
transform 1 0 11868 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0511_
timestamp 1632469394
transform 1 0 12972 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0509_
timestamp 1632469394
transform 1 0 12512 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1632469394
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_129
timestamp 1632469394
transform 1 0 12972 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1632469394
transform 1 0 12420 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _0516_
timestamp 1632469394
transform 1 0 13524 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1632469394
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0494_
timestamp 1632469394
transform 1 0 14352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1632469394
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1632469394
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1632469394
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0492_
timestamp 1632469394
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1632469394
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1632469394
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1632469394
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0761_
timestamp 1632469394
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0821_
timestamp 1632469394
transform 1 0 15824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0517_
timestamp 1632469394
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1632469394
transform 1 0 15640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1632469394
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1632469394
transform 1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1632469394
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1632469394
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1632469394
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1632469394
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1632469394
transform 1 0 17112 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0863_
timestamp 1632469394
transform 1 0 17112 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_14_173
timestamp 1632469394
transform 1 0 17020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 1632469394
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0877_
timestamp 1632469394
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 1632469394
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1632469394
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1632469394
transform 1 0 17572 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1632469394
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_189
timestamp 1632469394
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1632469394
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1632469394
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1632469394
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_196
timestamp 1632469394
transform 1 0 19136 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1632469394
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1632469394
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0521_
timestamp 1632469394
transform 1 0 19872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_200
timestamp 1632469394
transform 1 0 19504 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1632469394
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1632469394
transform 1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_208
timestamp 1632469394
transform 1 0 20240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_212
timestamp 1632469394
transform 1 0 20608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1632469394
transform -1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1632469394
transform -1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_216
timestamp 1632469394
transform 1 0 20976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1632469394
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1632469394
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1632469394
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0772_
timestamp 1632469394
transform 1 0 2116 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1632469394
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1632469394
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1632469394
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0787_
timestamp 1632469394
transform 1 0 4232 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0790_
timestamp 1632469394
transform 1 0 3128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1632469394
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1632469394
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1632469394
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0777_
timestamp 1632469394
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1632469394
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1632469394
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_84
timestamp 1632469394
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0778_
timestamp 1632469394
transform 1 0 7544 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1632469394
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1632469394
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1632469394
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_88
timestamp 1632469394
transform 1 0 9200 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1632469394
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1632469394
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0544_
timestamp 1632469394
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0716_
timestamp 1632469394
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1632469394
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1632469394
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 11776 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1632469394
transform 1 0 13248 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_136
timestamp 1632469394
transform 1 0 13616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1632469394
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_149
timestamp 1632469394
transform 1 0 14812 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0487_
timestamp 1632469394
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0561_
timestamp 1632469394
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1632469394
transform 1 0 15364 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1632469394
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1632469394
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1632469394
transform 1 0 16928 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1632469394
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0508_
timestamp 1632469394
transform 1 0 15456 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1632469394
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_180
timestamp 1632469394
transform 1 0 17664 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1632469394
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1632469394
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1632469394
transform 1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0528_
timestamp 1632469394
transform 1 0 18492 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_200
timestamp 1632469394
transform 1 0 19504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_207
timestamp 1632469394
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1632469394
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1632469394
transform -1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1632469394
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0524_
timestamp 1632469394
transform 1 0 19596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1632469394
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1632469394
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1632469394
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1632469394
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 2024 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1632469394
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_36
timestamp 1632469394
transform 1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_43
timestamp 1632469394
transform 1 0 5060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1632469394
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1632469394
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0758_
timestamp 1632469394
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_51
timestamp 1632469394
transform 1 0 5796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1632469394
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1632469394
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1632469394
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1632469394
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1632469394
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1632469394
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1632469394
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1632469394
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0762_
timestamp 1632469394
transform 1 0 7176 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_102
timestamp 1632469394
transform 1 0 10488 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1632469394
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1632469394
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0493_
timestamp 1632469394
transform 1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0532_
timestamp 1632469394
transform 1 0 10120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_116
timestamp 1632469394
transform 1 0 11776 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1632469394
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_1  _0513_
timestamp 1632469394
transform 1 0 12696 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0522_
timestamp 1632469394
transform 1 0 11224 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1632469394
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1632469394
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1632469394
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1632469394
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1632469394
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0489_
timestamp 1632469394
transform 1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1632469394
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1632469394
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0488_
timestamp 1632469394
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 15364 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 1632469394
transform 1 0 17112 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1632469394
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1632469394
transform 1 0 18308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1632469394
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1632469394
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1632469394
transform 1 0 18400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1632469394
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_210
timestamp 1632469394
transform 1 0 20424 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1632469394
transform -1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1632469394
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1632469394
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1632469394
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1632469394
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0760_
timestamp 1632469394
transform 1 0 2116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1632469394
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1632469394
transform 1 0 3864 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_37
timestamp 1632469394
transform 1 0 4508 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1632469394
transform 1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0771_
timestamp 1632469394
transform 1 0 3220 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1024_
timestamp 1632469394
transform 1 0 4876 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1632469394
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_63
timestamp 1632469394
transform 1 0 6900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1632469394
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0768_
timestamp 1632469394
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1632469394
transform 1 0 7636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_83
timestamp 1632469394
transform 1 0 8740 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0717_
timestamp 1632469394
transform 1 0 9108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp 1632469394
transform 1 0 7912 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1632469394
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1632469394
transform 1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1632469394
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1632469394
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1632469394
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1632469394
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _0514_
timestamp 1632469394
transform 1 0 12972 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0531_
timestamp 1632469394
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0533_
timestamp 1632469394
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1632469394
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_143
timestamp 1632469394
transform 1 0 14260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1632469394
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1632469394
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0495_
timestamp 1632469394
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1632469394
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1632469394
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1632469394
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0534_
timestamp 1632469394
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0967_
timestamp 1632469394
transform 1 0 15364 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1632469394
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1632469394
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0530_
timestamp 1632469394
transform 1 0 18032 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0540_
timestamp 1632469394
transform 1 0 19044 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_17_202
timestamp 1632469394
transform 1 0 19688 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1632469394
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_217
timestamp 1632469394
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1632469394
transform -1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0520_
timestamp 1632469394
transform 1 0 20240 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1632469394
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1632469394
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1632469394
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1632469394
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _0789_
timestamp 1632469394
transform 1 0 2668 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1632469394
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1632469394
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1632469394
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 1632469394
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1632469394
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1632469394
transform 1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1632469394
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1632469394
transform 1 0 6348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1632469394
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0755_
timestamp 1632469394
transform 1 0 5796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0767_
timestamp 1632469394
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1632469394
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1632469394
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _0763_
timestamp 1632469394
transform 1 0 7452 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 1632469394
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1632469394
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0620_
timestamp 1632469394
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1632469394
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1632469394
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_125
timestamp 1632469394
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0574_
timestamp 1632469394
transform 1 0 11500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0619_
timestamp 1632469394
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1632469394
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1632469394
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1632469394
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1632469394
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0647_
timestamp 1632469394
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0696_
timestamp 1632469394
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1632469394
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1632469394
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1632469394
transform 1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0535_
timestamp 1632469394
transform 1 0 17112 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1632469394
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1632469394
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_181
timestamp 1632469394
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1632469394
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1632469394
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1632469394
transform 1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1632469394
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1632469394
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_212
timestamp 1632469394
transform 1 0 20608 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1632469394
transform -1 0 21436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0542_
timestamp 1632469394
transform 1 0 20056 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1632469394
transform 1 0 19320 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1632469394
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1632469394
transform 1 0 1656 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1632469394
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1632469394
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1632469394
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1632469394
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0759_
timestamp 1632469394
transform 1 0 2668 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 1632469394
transform 1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1632469394
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_11
timestamp 1632469394
transform 1 0 2116 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1632469394
transform 1 0 3680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1632469394
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1632469394
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1632469394
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1632469394
transform 1 0 3312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0752_
timestamp 1632469394
transform 1 0 4692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1632469394
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1632469394
transform 1 0 4048 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1632469394
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_31
timestamp 1632469394
transform 1 0 3956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0753_
timestamp 1632469394
transform 1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_42
timestamp 1632469394
transform 1 0 4968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1632469394
transform 1 0 5336 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 1632469394
transform 1 0 5796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1632469394
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _0751_
timestamp 1632469394
transform 1 0 6624 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1632469394
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_59
timestamp 1632469394
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1632469394
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1632469394
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1632469394
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1632469394
transform 1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_65
timestamp 1632469394
transform 1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_75
timestamp 1632469394
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1632469394
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_67
timestamp 1632469394
transform 1 0 7268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1632469394
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1632469394
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1632469394
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0499_
timestamp 1632469394
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _0718_
timestamp 1632469394
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1632469394
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1632469394
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1632469394
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1632469394
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1632469394
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0711_
timestamp 1632469394
transform 1 0 10212 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  _0719_
timestamp 1632469394
transform 1 0 9200 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1632469394
transform 1 0 9936 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1632469394
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1632469394
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_126
timestamp 1632469394
transform 1 0 12696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1632469394
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_124
timestamp 1632469394
transform 1 0 12512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1632469394
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 1632469394
transform 1 0 12788 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1632469394
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1632469394
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1632469394
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1632469394
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1632469394
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1632469394
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0505_
timestamp 1632469394
transform 1 0 14720 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1632469394
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0695_
timestamp 1632469394
transform 1 0 13984 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1632469394
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1632469394
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1632469394
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1632469394
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1632469394
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0504_
timestamp 1632469394
transform 1 0 16652 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0507_
timestamp 1632469394
transform 1 0 15640 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0686_
timestamp 1632469394
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1632469394
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1632469394
transform 1 0 17572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0541_
timestamp 1632469394
transform 1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_175
timestamp 1632469394
transform 1 0 17204 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_182
timestamp 1632469394
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1632469394
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1632469394
transform 1 0 18400 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1632469394
transform 1 0 18584 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1632469394
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_184
timestamp 1632469394
transform 1 0 18032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1632469394
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_193
timestamp 1632469394
transform 1 0 18860 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1632469394
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _0543_
timestamp 1632469394
transform 1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1632469394
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1632469394
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1632469394
transform 1 0 20516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_214
timestamp 1632469394
transform 1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1632469394
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1632469394
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1632469394
transform -1 0 21436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1632469394
transform -1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1632469394
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1632469394
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1632469394
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0749_
timestamp 1632469394
transform 1 0 2116 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1632469394
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1632469394
transform 1 0 3496 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1632469394
transform 1 0 4232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1632469394
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1632469394
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0745_
timestamp 1632469394
transform 1 0 3128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 5060 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1632469394
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1632469394
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1632469394
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1632469394
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0750_
timestamp 1632469394
transform 1 0 6808 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1632469394
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1632469394
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1632469394
transform 1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1632469394
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_90
timestamp 1632469394
transform 1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1632469394
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0700_
timestamp 1632469394
transform 1 0 9660 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0710_
timestamp 1632469394
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1632469394
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1632469394
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1632469394
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1632469394
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0712_
timestamp 1632469394
transform 1 0 12788 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0715_
timestamp 1632469394
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1632469394
transform 1 0 13248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1632469394
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1632469394
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0689_
timestamp 1632469394
transform 1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0690_
timestamp 1632469394
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1632469394
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1632469394
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1632469394
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1020_
timestamp 1632469394
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1632469394
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1632469394
transform 1 0 18492 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _0545_
timestamp 1632469394
transform 1 0 17848 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0546_
timestamp 1632469394
transform 1 0 18860 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1632469394
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1632469394
transform 1 0 19872 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1632469394
transform 1 0 20700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_217
timestamp 1632469394
transform 1 0 21068 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1632469394
transform -1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0552_
timestamp 1632469394
transform 1 0 19964 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1632469394
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1632469394
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1632469394
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1632469394
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0746_
timestamp 1632469394
transform 1 0 2300 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1632469394
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1632469394
transform 1 0 4048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1632469394
transform 1 0 4784 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1632469394
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _0739_
timestamp 1632469394
transform 1 0 4876 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1632469394
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1632469394
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1632469394
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1632469394
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _0737_
timestamp 1632469394
transform 1 0 6808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1632469394
transform 1 0 5704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1632469394
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1632469394
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1632469394
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1632469394
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0697_
timestamp 1632469394
transform 1 0 9016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_109
timestamp 1632469394
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_89
timestamp 1632469394
transform 1 0 9292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1632469394
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0698_
timestamp 1632469394
transform 1 0 9660 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0709_
timestamp 1632469394
transform 1 0 10580 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1632469394
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1632469394
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0728_
timestamp 1632469394
transform 1 0 12880 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0729_
timestamp 1632469394
transform 1 0 11776 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1632469394
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1632469394
transform 1 0 14720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1632469394
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1632469394
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0694_
timestamp 1632469394
transform 1 0 14076 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_155
timestamp 1632469394
transform 1 0 15364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_163
timestamp 1632469394
transform 1 0 16100 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_169
timestamp 1632469394
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0684_
timestamp 1632469394
transform 1 0 17020 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1632469394
transform 1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1632469394
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_181
timestamp 1632469394
transform 1 0 17756 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1632469394
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1632469394
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0683_
timestamp 1632469394
transform 1 0 17848 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1632469394
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1632469394
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_214
timestamp 1632469394
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1632469394
transform -1 0 21436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0536_
timestamp 1632469394
transform 1 0 20332 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0539_
timestamp 1632469394
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1632469394
transform 1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1632469394
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1632469394
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1632469394
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0733_
timestamp 1632469394
transform 1 0 2668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1632469394
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_25
timestamp 1632469394
transform 1 0 3404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_33
timestamp 1632469394
transform 1 0 4140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_40
timestamp 1632469394
transform 1 0 4784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0721_
timestamp 1632469394
transform 1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1632469394
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1632469394
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1632469394
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0736_
timestamp 1632469394
transform 1 0 6900 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0741_
timestamp 1632469394
transform 1 0 5336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_72
timestamp 1632469394
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_84
timestamp 1632469394
transform 1 0 8832 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1632469394
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1632469394
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1632469394
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1632469394
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1632469394
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1632469394
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_126
timestamp 1632469394
transform 1 0 12696 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1632469394
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_2  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1632469394
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_151
timestamp 1632469394
transform 1 0 14996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1632469394
transform 1 0 13432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _0704_
timestamp 1632469394
transform 1 0 14076 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1632469394
transform 1 0 15364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1632469394
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1632469394
transform 1 0 16928 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1632469394
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1632469394
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0726_
timestamp 1632469394
transform 1 0 15456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1632469394
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_185
timestamp 1632469394
transform 1 0 18124 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_193
timestamp 1632469394
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1632469394
transform 1 0 17848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1632469394
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1632469394
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_211
timestamp 1632469394
transform 1 0 20516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_217
timestamp 1632469394
transform 1 0 21068 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1632469394
transform -1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 1632469394
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1632469394
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1632469394
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0735_
timestamp 1632469394
transform 1 0 2668 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1632469394
transform 1 0 1380 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1632469394
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1632469394
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1632469394
transform 1 0 4968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1632469394
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1632469394
transform 1 0 4140 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1632469394
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1632469394
transform 1 0 6808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1632469394
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1632469394
transform 1 0 5336 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_72
timestamp 1632469394
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1632469394
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _0503_
timestamp 1632469394
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0723_
timestamp 1632469394
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1632469394
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1632469394
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0707_
timestamp 1632469394
transform 1 0 9844 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0714_
timestamp 1632469394
transform 1 0 10856 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_113
timestamp 1632469394
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1632469394
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1632469394
transform 1 0 11868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0725_
timestamp 1632469394
transform 1 0 12880 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1632469394
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1632469394
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1632469394
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_147
timestamp 1632469394
transform 1 0 14628 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1632469394
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1632469394
transform 1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_162
timestamp 1632469394
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1632469394
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1632469394
transform 1 0 16928 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0671_
timestamp 1632469394
transform 1 0 15364 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_175
timestamp 1632469394
transform 1 0 17204 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_183
timestamp 1632469394
transform 1 0 17940 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1632469394
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1632469394
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1632469394
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0666_
timestamp 1632469394
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_200
timestamp 1632469394
transform 1 0 19504 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_214
timestamp 1632469394
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1632469394
transform -1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1632469394
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1632469394
transform 1 0 19872 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_25_14
timestamp 1632469394
transform 1 0 2392 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_20
timestamp 1632469394
transform 1 0 2944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1632469394
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1632469394
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0788_
timestamp 1632469394
transform 1 0 3036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0983_
timestamp 1632469394
transform 1 0 1564 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_29
timestamp 1632469394
transform 1 0 3772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_36
timestamp 1632469394
transform 1 0 4416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0740_
timestamp 1632469394
transform 1 0 4784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1632469394
transform 1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1632469394
transform 1 0 5152 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1632469394
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1632469394
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1632469394
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1632469394
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1632469394
transform 1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 1632469394
transform 1 0 6716 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1632469394
transform 1 0 7544 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1632469394
transform 1 0 8648 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 1632469394
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0706_
timestamp 1632469394
transform 1 0 9752 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1632469394
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1632469394
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1632469394
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1632469394
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1632469394
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1632469394
transform 1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0705_
timestamp 1632469394
transform 1 0 11776 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_25_138
timestamp 1632469394
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_151
timestamp 1632469394
transform 1 0 14996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0691_
timestamp 1632469394
transform 1 0 14352 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0727_
timestamp 1632469394
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1632469394
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1632469394
transform 1 0 16928 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1632469394
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1632469394
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0680_
timestamp 1632469394
transform 1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_185
timestamp 1632469394
transform 1 0 18124 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1632469394
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1632469394
transform 1 0 17296 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1632469394
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_199
timestamp 1632469394
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_211
timestamp 1632469394
transform 1 0 20516 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1632469394
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1632469394
transform -1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0537_
timestamp 1632469394
transform 1 0 19780 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1632469394
transform 1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 1632469394
transform 1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1632469394
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1632469394
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1632469394
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1632469394
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1632469394
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1632469394
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1632469394
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_14
timestamp 1632469394
transform 1 0 2392 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_10
timestamp 1632469394
transform 1 0 2024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1632469394
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_18
timestamp 1632469394
transform 1 0 2760 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1632469394
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1632469394
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0575_
timestamp 1632469394
transform 1 0 3588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1632469394
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_26
timestamp 1632469394
transform 1 0 3496 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1632469394
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1632469394
transform 1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_33
timestamp 1632469394
transform 1 0 4140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1632469394
transform 1 0 4692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1632469394
transform 1 0 4048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0581_
timestamp 1632469394
transform 1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0579_
timestamp 1632469394
transform 1 0 5060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_41
timestamp 1632469394
transform 1 0 4876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1632469394
transform 1 0 5888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1632469394
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_51
timestamp 1632469394
transform 1 0 5796 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1632469394
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0582_
timestamp 1632469394
transform 1 0 6808 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0565_
timestamp 1632469394
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1632469394
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_60
timestamp 1632469394
transform 1 0 6624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1632469394
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1632469394
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_55
timestamp 1632469394
transform 1 0 6164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  _0583_
timestamp 1632469394
transform 1 0 6992 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_26_71
timestamp 1632469394
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1632469394
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1632469394
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_71
timestamp 1632469394
transform 1 0 7636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_79
timestamp 1632469394
transform 1 0 8372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_86
timestamp 1632469394
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1632469394
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0560_
timestamp 1632469394
transform 1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1632469394
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1632469394
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1632469394
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1632469394
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1632469394
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1632469394
transform 1 0 10672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 1632469394
transform 1 0 9752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1632469394
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1632469394
transform 1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1632469394
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1632469394
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1632469394
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_116
timestamp 1632469394
transform 1 0 11776 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1632469394
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_117
timestamp 1632469394
transform 1 0 11868 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1632469394
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1632469394
transform 1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0562_
timestamp 1632469394
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1632469394
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1632469394
transform 1 0 12604 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1632469394
transform 1 0 12880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_131
timestamp 1632469394
transform 1 0 13156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1632469394
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1632469394
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_148
timestamp 1632469394
transform 1 0 14720 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_148
timestamp 1632469394
transform 1 0 14720 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1632469394
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _0678_
timestamp 1632469394
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1632469394
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 1632469394
transform 1 0 13892 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_1  _0681_
timestamp 1632469394
transform 1 0 15548 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0506_
timestamp 1632469394
transform 1 0 15364 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1632469394
transform 1 0 15272 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_156
timestamp 1632469394
transform 1 0 15456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1632469394
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1632469394
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1632469394
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_164
timestamp 1632469394
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1632469394
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _0556_
timestamp 1632469394
transform 1 0 17112 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1632469394
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1632469394
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1632469394
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0668_
timestamp 1632469394
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_181
timestamp 1632469394
transform 1 0 17756 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1632469394
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0549_
timestamp 1632469394
transform 1 0 18216 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1632469394
transform 1 0 18400 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_27_187
timestamp 1632469394
transform 1 0 18308 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1632469394
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1632469394
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1632469394
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1632469394
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1632469394
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0551_
timestamp 1632469394
transform 1 0 19320 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1632469394
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_197
timestamp 1632469394
transform 1 0 19228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1632469394
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_1  _0554_
timestamp 1632469394
transform 1 0 20240 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1632469394
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_216
timestamp 1632469394
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_208
timestamp 1632469394
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1632469394
transform -1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1632469394
transform -1 0 21436 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_11
timestamp 1632469394
transform 1 0 2116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_17
timestamp 1632469394
transform 1 0 2668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1632469394
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1632469394
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0572_
timestamp 1632469394
transform 1 0 2760 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1632469394
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1632469394
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1632469394
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_42
timestamp 1632469394
transform 1 0 4968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1632469394
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0580_
timestamp 1632469394
transform 1 0 5060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1632469394
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1632469394
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1632469394
transform 1 0 6624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0566_
timestamp 1632469394
transform 1 0 5980 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1632469394
transform 1 0 6992 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1632469394
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_73
timestamp 1632469394
transform 1 0 7820 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1632469394
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1632469394
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0563_
timestamp 1632469394
transform 1 0 7912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _0568_
timestamp 1632469394
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_28_103
timestamp 1632469394
transform 1 0 10580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_92
timestamp 1632469394
transform 1 0 9568 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _0621_
timestamp 1632469394
transform 1 0 9936 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1632469394
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_121
timestamp 1632469394
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_128
timestamp 1632469394
transform 1 0 12880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1632469394
transform 1 0 11960 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1632469394
transform 1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1632469394
transform 1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_132
timestamp 1632469394
transform 1 0 13248 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1632469394
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1632469394
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1632469394
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1632469394
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0677_
timestamp 1632469394
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 1632469394
transform 1 0 13340 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1632469394
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1632469394
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1632469394
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1632469394
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _0664_
timestamp 1632469394
transform 1 0 15640 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1632469394
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1632469394
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1632469394
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _0557_
timestamp 1632469394
transform 1 0 18124 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0559_
timestamp 1632469394
transform 1 0 17296 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1632469394
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1632469394
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_214
timestamp 1632469394
transform 1 0 20792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1632469394
transform -1 0 21436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0553_
timestamp 1632469394
transform 1 0 20516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0564_
timestamp 1632469394
transform 1 0 19412 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_17
timestamp 1632469394
transform 1 0 2668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1632469394
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_8
timestamp 1632469394
transform 1 0 1840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1632469394
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0567_
timestamp 1632469394
transform 1 0 3036 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0570_
timestamp 1632469394
transform 1 0 2208 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1632469394
transform 1 0 1472 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1632469394
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_35
timestamp 1632469394
transform 1 0 4324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1632469394
transform 1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1632469394
transform 1 0 4048 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1632469394
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_65
timestamp 1632469394
transform 1 0 7084 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1632469394
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0591_
timestamp 1632469394
transform 1 0 5244 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0612_
timestamp 1632469394
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1632469394
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0569_
timestamp 1632469394
transform 1 0 7820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1632469394
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1632469394
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1632469394
transform 1 0 10488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1632469394
transform 1 0 9292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1632469394
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_120
timestamp 1632469394
transform 1 0 12144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_131
timestamp 1632469394
transform 1 0 13156 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1632469394
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0618_
timestamp 1632469394
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0634_
timestamp 1632469394
transform 1 0 12512 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1632469394
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_142
timestamp 1632469394
transform 1 0 14168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_146
timestamp 1632469394
transform 1 0 14536 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1632469394
transform 1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1632469394
transform 1 0 14260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_154
timestamp 1632469394
transform 1 0 15272 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1632469394
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1632469394
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1632469394
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1632469394
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0654_
timestamp 1632469394
transform 1 0 17112 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0663_
timestamp 1632469394
transform 1 0 15364 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1632469394
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1632469394
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_188
timestamp 1632469394
transform 1 0 18400 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_194
timestamp 1632469394
transform 1 0 18952 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1632469394
transform 1 0 18124 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1632469394
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1632469394
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_211
timestamp 1632469394
transform 1 0 20516 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1632469394
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1632469394
transform -1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0555_
timestamp 1632469394
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1632469394
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1632469394
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1632469394
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1632469394
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1632469394
transform 1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1632469394
transform 1 0 1564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1632469394
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1632469394
transform 1 0 4048 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1632469394
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1632469394
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1632469394
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1632469394
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1632469394
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1632469394
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1632469394
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0613_
timestamp 1632469394
transform 1 0 5336 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 1632469394
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1632469394
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_66
timestamp 1632469394
transform 1 0 7176 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_74
timestamp 1632469394
transform 1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1632469394
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1632469394
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1632469394
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1632469394
transform 1 0 9016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1632469394
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_104
timestamp 1632469394
transform 1 0 10672 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_89
timestamp 1632469394
transform 1 0 9292 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 1632469394
transform 1 0 9844 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_110
timestamp 1632469394
transform 1 0 11224 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_119
timestamp 1632469394
transform 1 0 12052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_123
timestamp 1632469394
transform 1 0 12420 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _0615_
timestamp 1632469394
transform 1 0 11316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 1632469394
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1632469394
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1632469394
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1632469394
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1632469394
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_1  _0672_
timestamp 1632469394
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1632469394
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1632469394
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0657_
timestamp 1632469394
transform 1 0 16284 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0676_
timestamp 1632469394
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_185
timestamp 1632469394
transform 1 0 18124 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1632469394
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1632469394
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1632469394
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1632469394
transform 1 0 17296 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1632469394
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_210
timestamp 1632469394
transform 1 0 20424 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1632469394
transform -1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 1632469394
transform 1 0 19596 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_16
timestamp 1632469394
transform 1 0 2576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1632469394
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1632469394
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0585_
timestamp 1632469394
transform 1 0 2116 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0596_
timestamp 1632469394
transform 1 0 2944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1632469394
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_28
timestamp 1632469394
transform 1 0 3680 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_38
timestamp 1632469394
transform 1 0 4600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1632469394
transform 1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0598_
timestamp 1632469394
transform 1 0 4048 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 1632469394
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1632469394
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1632469394
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1632469394
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632469394
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1632469394
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1632469394
transform 1 0 7912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_81
timestamp 1632469394
transform 1 0 8556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_85
timestamp 1632469394
transform 1 0 8924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1632469394
transform 1 0 8280 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0609_
timestamp 1632469394
transform 1 0 9016 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1632469394
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_103
timestamp 1632469394
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_92
timestamp 1632469394
transform 1 0 9568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _0622_
timestamp 1632469394
transform 1 0 9936 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1632469394
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1632469394
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1632469394
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1632469394
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1632469394
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1632469394
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0631_
timestamp 1632469394
transform 1 0 11960 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_31_132
timestamp 1632469394
transform 1 0 13248 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1632469394
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1632469394
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1632469394
transform 1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _0675_
timestamp 1632469394
transform 1 0 13800 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_31_156
timestamp 1632469394
transform 1 0 15456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1632469394
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1632469394
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1632469394
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1632469394
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0673_
timestamp 1632469394
transform 1 0 15548 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1632469394
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_185
timestamp 1632469394
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1632469394
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _0652_
timestamp 1632469394
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1632469394
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1632469394
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1632469394
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_214
timestamp 1632469394
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1632469394
transform -1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1632469394
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1632469394
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_13
timestamp 1632469394
transform 1 0 2300 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1632469394
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0595_
timestamp 1632469394
transform 1 0 2852 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1632469394
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1632469394
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_38
timestamp 1632469394
transform 1 0 4600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1632469394
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 1632469394
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_46
timestamp 1632469394
transform 1 0 5336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1632469394
transform 1 0 5888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_60
timestamp 1632469394
transform 1 0 6624 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0604_
timestamp 1632469394
transform 1 0 6992 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0611_
timestamp 1632469394
transform 1 0 5428 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1632469394
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_73
timestamp 1632469394
transform 1 0 7820 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1632469394
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1632469394
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1632469394
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1632469394
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_100
timestamp 1632469394
transform 1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1632469394
transform 1 0 11040 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1632469394
transform 1 0 9476 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1632469394
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_115
timestamp 1632469394
transform 1 0 11684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1632469394
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_128
timestamp 1632469394
transform 1 0 12880 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1632469394
transform 1 0 11408 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0674_
timestamp 1632469394
transform 1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1632469394
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1632469394
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1632469394
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1632469394
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1632469394
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1632469394
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1632469394
transform 1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1632469394
transform 1 0 15548 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1632469394
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1632469394
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1632469394
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1632469394
transform 1 0 15640 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1632469394
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1632469394
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1632469394
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1632469394
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1632469394
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1632469394
transform 1 0 18400 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1632469394
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1632469394
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1632469394
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1632469394
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1632469394
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1632469394
transform -1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1632469394
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1632469394
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1632469394
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1632469394
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1632469394
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1632469394
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1632469394
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_7
timestamp 1632469394
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1632469394
transform 1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1632469394
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1632469394
transform 1 0 2116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1632469394
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0586_
timestamp 1632469394
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1632469394
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1632469394
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0587_
timestamp 1632469394
transform 1 0 3680 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1632469394
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1632469394
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1632469394
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_23
timestamp 1632469394
transform 1 0 3220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1632469394
transform 1 0 4600 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_38
timestamp 1632469394
transform 1 0 4600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1632469394
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1632469394
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1632469394
transform 1 0 4968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0610_
timestamp 1632469394
transform 1 0 5244 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0590_
timestamp 1632469394
transform 1 0 5704 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_46
timestamp 1632469394
transform 1 0 5336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0601_
timestamp 1632469394
transform 1 0 6348 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1632469394
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1632469394
transform 1 0 6348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1632469394
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1632469394
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_65
timestamp 1632469394
transform 1 0 7084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_64
timestamp 1632469394
transform 1 0 6992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_70
timestamp 1632469394
transform 1 0 7544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_78
timestamp 1632469394
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1632469394
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1632469394
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1632469394
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_1  _0593_
timestamp 1632469394
transform 1 0 7452 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_1  _0594_
timestamp 1632469394
transform 1 0 7636 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0605_
timestamp 1632469394
transform 1 0 8648 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1632469394
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1632469394
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1632469394
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_105
timestamp 1632469394
transform 1 0 10764 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1632469394
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0607_
timestamp 1632469394
transform 1 0 9660 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0624_
timestamp 1632469394
transform 1 0 10580 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0625_
timestamp 1632469394
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1632469394
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_1  _0636_
timestamp 1632469394
transform 1 0 11592 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0635_
timestamp 1632469394
transform 1 0 11408 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1632469394
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_111
timestamp 1632469394
transform 1 0 11316 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1632469394
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _0646_
timestamp 1632469394
transform 1 0 12880 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0645_
timestamp 1632469394
transform 1 0 12696 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1632469394
transform 1 0 12788 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_121
timestamp 1632469394
transform 1 0 12236 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1632469394
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_121
timestamp 1632469394
transform 1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1632469394
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_137
timestamp 1632469394
transform 1 0 13708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1632469394
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1632469394
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1632469394
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1632469394
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0661_
timestamp 1632469394
transform 1 0 14536 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp 1632469394
transform 1 0 14352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1632469394
transform 1 0 13800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1632469394
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1632469394
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1632469394
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1632469394
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1632469394
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1632469394
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0644_
timestamp 1632469394
transform 1 0 15548 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0648_
timestamp 1632469394
transform 1 0 16100 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_1  _0649_
timestamp 1632469394
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1022_
timestamp 1632469394
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0641_
timestamp 1632469394
transform 1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_176
timestamp 1632469394
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0651_
timestamp 1632469394
transform 1 0 18584 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1632469394
transform 1 0 18492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1632469394
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1632469394
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1632469394
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1632469394
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_195
timestamp 1632469394
transform 1 0 19044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1632469394
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1632469394
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1632469394
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1632469394
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1632469394
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1632469394
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1632469394
transform 1 0 20424 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_209
timestamp 1632469394
transform 1 0 20332 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1632469394
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1632469394
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1632469394
transform -1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1632469394
transform -1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_217
timestamp 1632469394
transform 1 0 21068 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1632469394
transform 1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_19
timestamp 1632469394
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1632469394
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1632469394
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1632469394
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1632469394
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1632469394
transform 1 0 3588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_38
timestamp 1632469394
transform 1 0 4600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0603_
timestamp 1632469394
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp 1632469394
transform 1 0 3772 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1632469394
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_64
timestamp 1632469394
transform 1 0 6992 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1632469394
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _0592_
timestamp 1632469394
transform 1 0 6348 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1632469394
transform 1 0 7728 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_83
timestamp 1632469394
transform 1 0 8740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1632469394
transform 1 0 7912 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1632469394
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_93
timestamp 1632469394
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0626_
timestamp 1632469394
transform 1 0 10028 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1632469394
transform 1 0 9292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1632469394
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_117
timestamp 1632469394
transform 1 0 11868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1632469394
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1632469394
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _0630_
timestamp 1632469394
transform 1 0 12236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp 1632469394
transform 1 0 12972 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1632469394
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1632469394
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1632469394
transform 1 0 14444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0629_
timestamp 1632469394
transform 1 0 14168 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0658_
timestamp 1632469394
transform 1 0 14812 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_156
timestamp 1632469394
transform 1 0 15456 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1632469394
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1632469394
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_174
timestamp 1632469394
transform 1 0 17112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1632469394
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1632469394
transform 1 0 16744 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1632469394
transform 1 0 15824 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1632469394
transform 1 0 18032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1632469394
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1632469394
transform 1 0 18400 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0639_
timestamp 1632469394
transform 1 0 17480 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1632469394
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1632469394
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1632469394
transform -1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1632469394
transform 1 0 19228 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1632469394
transform 1 0 19872 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_36_11
timestamp 1632469394
transform 1 0 2116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_19
timestamp 1632469394
transform 1 0 2852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1632469394
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1632469394
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1632469394
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1632469394
transform 1 0 2944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1632469394
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1632469394
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_43
timestamp 1632469394
transform 1 0 5060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1632469394
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1632469394
transform 1 0 4140 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_36_47
timestamp 1632469394
transform 1 0 5428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_52
timestamp 1632469394
transform 1 0 5888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_64
timestamp 1632469394
transform 1 0 6992 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1632469394
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0602_
timestamp 1632469394
transform 1 0 6348 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1632469394
transform 1 0 5520 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_70
timestamp 1632469394
transform 1 0 7544 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_75
timestamp 1632469394
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1632469394
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1632469394
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1632469394
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1632469394
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_101
timestamp 1632469394
transform 1 0 10396 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1632469394
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1632469394
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0606_
timestamp 1632469394
transform 1 0 10764 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1632469394
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1632469394
transform 1 0 9292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1632469394
transform 1 0 12420 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1632469394
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1632469394
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1632469394
transform 1 0 11500 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1632469394
transform 1 0 12788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1632469394
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1632469394
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1632469394
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1632469394
transform 1 0 14812 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1632469394
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_159
timestamp 1632469394
transform 1 0 15732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_167
timestamp 1632469394
transform 1 0 16468 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1632469394
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1632469394
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1632469394
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_177
timestamp 1632469394
transform 1 0 17388 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_185
timestamp 1632469394
transform 1 0 18124 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1632469394
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1632469394
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1632469394
transform 1 0 18400 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_200
timestamp 1632469394
transform 1 0 19504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1632469394
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1632469394
transform -1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1632469394
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1632469394
transform 1 0 19872 0 1 21760
box -38 -48 958 592
<< labels >>
rlabel metal2 s 14738 23911 14794 24711 6 A[0]
port 0 nsew signal input
rlabel metal3 s 21767 16600 22567 16720 6 A[10]
port 1 nsew signal input
rlabel metal3 s 21767 5176 22567 5296 6 A[11]
port 2 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 A[12]
port 3 nsew signal input
rlabel metal3 s 21767 12248 22567 12368 6 A[13]
port 4 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 A[14]
port 5 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 A[15]
port 6 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 A[16]
port 7 nsew signal input
rlabel metal2 s 19522 23911 19578 24711 6 A[17]
port 8 nsew signal input
rlabel metal2 s 5906 23911 5962 24711 6 A[18]
port 9 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 A[19]
port 10 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 A[1]
port 11 nsew signal input
rlabel metal3 s 21767 18504 22567 18624 6 A[20]
port 12 nsew signal input
rlabel metal2 s 21914 23911 21970 24711 6 A[21]
port 13 nsew signal input
rlabel metal3 s 0 824 800 944 6 A[22]
port 14 nsew signal input
rlabel metal3 s 21767 17688 22567 17808 6 A[23]
port 15 nsew signal input
rlabel metal3 s 21767 7080 22567 7200 6 A[24]
port 16 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 A[25]
port 17 nsew signal input
rlabel metal2 s 16578 23911 16634 24711 6 A[26]
port 18 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 A[27]
port 19 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 A[28]
port 20 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 A[29]
port 21 nsew signal input
rlabel metal3 s 21767 14968 22567 15088 6 A[2]
port 22 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 A[30]
port 23 nsew signal input
rlabel metal2 s 9954 23911 10010 24711 6 A[31]
port 24 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 A[3]
port 25 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 A[4]
port 26 nsew signal input
rlabel metal2 s 20258 23911 20314 24711 6 A[5]
port 27 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 A[6]
port 28 nsew signal input
rlabel metal3 s 21767 13064 22567 13184 6 A[7]
port 29 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 A[8]
port 30 nsew signal input
rlabel metal3 s 21767 22040 22567 22160 6 A[9]
port 31 nsew signal input
rlabel metal3 s 21767 7896 22567 8016 6 B[0]
port 32 nsew signal input
rlabel metal2 s 4066 23911 4122 24711 6 B[10]
port 33 nsew signal input
rlabel metal3 s 21767 23672 22567 23792 6 B[11]
port 34 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 B[12]
port 35 nsew signal input
rlabel metal3 s 21767 3544 22567 3664 6 B[13]
port 36 nsew signal input
rlabel metal2 s 10690 23911 10746 24711 6 B[14]
port 37 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 B[15]
port 38 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 B[16]
port 39 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 B[17]
port 40 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 B[18]
port 41 nsew signal input
rlabel metal2 s 13082 23911 13138 24711 6 B[19]
port 42 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 B[1]
port 43 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 B[20]
port 44 nsew signal input
rlabel metal2 s 5170 23911 5226 24711 6 B[21]
port 45 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 B[22]
port 46 nsew signal input
rlabel metal2 s 570 0 626 800 6 B[23]
port 47 nsew signal input
rlabel metal2 s 16026 23911 16082 24711 6 B[24]
port 48 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 B[25]
port 49 nsew signal input
rlabel metal2 s 21362 23911 21418 24711 6 B[26]
port 50 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 B[27]
port 51 nsew signal input
rlabel metal2 s 8298 23911 8354 24711 6 B[28]
port 52 nsew signal input
rlabel metal2 s 3514 23911 3570 24711 6 B[29]
port 53 nsew signal input
rlabel metal2 s 7562 23911 7618 24711 6 B[2]
port 54 nsew signal input
rlabel metal2 s 12346 23911 12402 24711 6 B[30]
port 55 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 B[31]
port 56 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 B[3]
port 57 nsew signal input
rlabel metal2 s 22466 23911 22522 24711 6 B[4]
port 58 nsew signal input
rlabel metal2 s 1674 23911 1730 24711 6 B[5]
port 59 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 B[6]
port 60 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 B[7]
port 61 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 B[8]
port 62 nsew signal input
rlabel metal2 s 13634 23911 13690 24711 6 B[9]
port 63 nsew signal input
rlabel metal3 s 21767 20136 22567 20256 6 Enable
port 64 nsew signal input
rlabel metal2 s 18970 23911 19026 24711 6 Result[0]
port 65 nsew signal tristate
rlabel metal2 s 4618 23911 4674 24711 6 Result[10]
port 66 nsew signal tristate
rlabel metal2 s 9402 23911 9458 24711 6 Result[11]
port 67 nsew signal tristate
rlabel metal2 s 11242 23911 11298 24711 6 Result[12]
port 68 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 Result[13]
port 69 nsew signal tristate
rlabel metal2 s 7010 23911 7066 24711 6 Result[14]
port 70 nsew signal tristate
rlabel metal3 s 21767 4360 22567 4480 6 Result[15]
port 71 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 Result[16]
port 72 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 Result[17]
port 73 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 Result[18]
port 74 nsew signal tristate
rlabel metal3 s 21767 5992 22567 6112 6 Result[19]
port 75 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 Result[1]
port 76 nsew signal tristate
rlabel metal3 s 21767 1640 22567 1760 6 Result[20]
port 77 nsew signal tristate
rlabel metal3 s 0 5176 800 5296 6 Result[21]
port 78 nsew signal tristate
rlabel metal2 s 8850 0 8906 800 6 Result[22]
port 79 nsew signal tristate
rlabel metal3 s 21767 10616 22567 10736 6 Result[23]
port 80 nsew signal tristate
rlabel metal3 s 21767 22856 22567 22976 6 Result[24]
port 81 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 Result[25]
port 82 nsew signal tristate
rlabel metal3 s 21767 8 22567 128 6 Result[26]
port 83 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 Result[27]
port 84 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 Result[28]
port 85 nsew signal tristate
rlabel metal2 s 11794 23911 11850 24711 6 Result[29]
port 86 nsew signal tristate
rlabel metal2 s 14922 0 14978 800 6 Result[2]
port 87 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 Result[30]
port 88 nsew signal tristate
rlabel metal3 s 0 10344 800 10464 6 Result[31]
port 89 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 Result[32]
port 90 nsew signal tristate
rlabel metal3 s 21767 15784 22567 15904 6 Result[33]
port 91 nsew signal tristate
rlabel metal3 s 21767 8712 22567 8832 6 Result[34]
port 92 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 Result[35]
port 93 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 Result[36]
port 94 nsew signal tristate
rlabel metal3 s 21767 2456 22567 2576 6 Result[37]
port 95 nsew signal tristate
rlabel metal3 s 0 1640 800 1760 6 Result[38]
port 96 nsew signal tristate
rlabel metal3 s 21767 11432 22567 11552 6 Result[39]
port 97 nsew signal tristate
rlabel metal3 s 21767 19320 22567 19440 6 Result[3]
port 98 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 Result[40]
port 99 nsew signal tristate
rlabel metal3 s 21767 21224 22567 21344 6 Result[41]
port 100 nsew signal tristate
rlabel metal2 s 570 23911 626 24711 6 Result[42]
port 101 nsew signal tristate
rlabel metal3 s 0 13064 800 13184 6 Result[43]
port 102 nsew signal tristate
rlabel metal2 s 10690 0 10746 800 6 Result[44]
port 103 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 Result[45]
port 104 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 Result[46]
port 105 nsew signal tristate
rlabel metal2 s 2226 23911 2282 24711 6 Result[47]
port 106 nsew signal tristate
rlabel metal2 s 8850 23911 8906 24711 6 Result[48]
port 107 nsew signal tristate
rlabel metal2 s 15474 23911 15530 24711 6 Result[49]
port 108 nsew signal tristate
rlabel metal3 s 0 22856 800 22976 6 Result[4]
port 109 nsew signal tristate
rlabel metal3 s 0 11432 800 11552 6 Result[50]
port 110 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 Result[51]
port 111 nsew signal tristate
rlabel metal2 s 18418 23911 18474 24711 6 Result[52]
port 112 nsew signal tristate
rlabel metal2 s 14186 23911 14242 24711 6 Result[53]
port 113 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 Result[54]
port 114 nsew signal tristate
rlabel metal2 s 20810 23911 20866 24711 6 Result[55]
port 115 nsew signal tristate
rlabel metal3 s 21767 824 22567 944 6 Result[56]
port 116 nsew signal tristate
rlabel metal2 s 1122 23911 1178 24711 6 Result[57]
port 117 nsew signal tristate
rlabel metal3 s 0 8712 800 8832 6 Result[58]
port 118 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 Result[59]
port 119 nsew signal tristate
rlabel metal2 s 7010 0 7066 800 6 Result[5]
port 120 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 Result[60]
port 121 nsew signal tristate
rlabel metal3 s 21767 14152 22567 14272 6 Result[61]
port 122 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 Result[62]
port 123 nsew signal tristate
rlabel metal2 s 17866 23911 17922 24711 6 Result[63]
port 124 nsew signal tristate
rlabel metal2 s 17130 23911 17186 24711 6 Result[6]
port 125 nsew signal tristate
rlabel metal2 s 2778 23911 2834 24711 6 Result[7]
port 126 nsew signal tristate
rlabel metal2 s 6458 23911 6514 24711 6 Result[8]
port 127 nsew signal tristate
rlabel metal2 s 13634 0 13690 800 6 Result[9]
port 128 nsew signal tristate
rlabel metal5 s 1104 8677 21436 8997 6 VGND
port 129 nsew ground input
rlabel metal5 s 1104 15386 21436 15706 6 VGND
port 129 nsew ground input
rlabel metal4 s 7721 2128 8041 22352 6 VGND
port 129 nsew ground input
rlabel metal4 s 14498 2128 14818 22352 6 VGND
port 129 nsew ground input
rlabel metal5 s 1104 5323 21436 5643 6 VPWR
port 130 nsew power input
rlabel metal5 s 1104 12032 21436 12352 6 VPWR
port 130 nsew power input
rlabel metal5 s 1104 18741 21436 19061 6 VPWR
port 130 nsew power input
rlabel metal4 s 4333 2128 4653 22352 6 VPWR
port 130 nsew power input
rlabel metal4 s 11110 2128 11430 22352 6 VPWR
port 130 nsew power input
rlabel metal4 s 17887 2128 18207 22352 6 VPWR
port 130 nsew power input
rlabel metal3 s 0 7896 800 8016 6 opcode[0]
port 131 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 opcode[1]
port 132 nsew signal input
rlabel metal3 s 21767 9528 22567 9648 6 opcode[2]
port 133 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 22567 24711
<< end >>
