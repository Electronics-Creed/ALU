VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu32
  CLASS BLOCK ;
  FOREIGN alu32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 112.835 BY 123.555 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 119.555 73.970 123.555 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 83.000 112.835 83.600 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 25.880 112.835 26.480 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 61.240 112.835 61.840 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 119.555 97.890 123.555 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 119.555 29.810 123.555 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 92.520 112.835 93.120 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 119.555 109.850 123.555 ;
    END
  END A[21]
  PIN A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END A[22]
  PIN A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 88.440 112.835 89.040 ;
    END
  END A[23]
  PIN A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 35.400 112.835 36.000 ;
    END
  END A[24]
  PIN A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END A[25]
  PIN A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 119.555 83.170 123.555 ;
    END
  END A[26]
  PIN A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END A[27]
  PIN A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END A[28]
  PIN A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END A[29]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 74.840 112.835 75.440 ;
    END
  END A[2]
  PIN A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END A[30]
  PIN A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 119.555 50.050 123.555 ;
    END
  END A[31]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 119.555 101.570 123.555 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 65.320 112.835 65.920 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 110.200 112.835 110.800 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 39.480 112.835 40.080 ;
    END
  END B[0]
  PIN B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 119.555 20.610 123.555 ;
    END
  END B[10]
  PIN B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 118.360 112.835 118.960 ;
    END
  END B[11]
  PIN B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END B[12]
  PIN B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 17.720 112.835 18.320 ;
    END
  END B[13]
  PIN B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 119.555 53.730 123.555 ;
    END
  END B[14]
  PIN B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END B[15]
  PIN B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END B[16]
  PIN B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END B[17]
  PIN B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END B[18]
  PIN B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 119.555 65.690 123.555 ;
    END
  END B[19]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END B[1]
  PIN B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END B[20]
  PIN B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 119.555 26.130 123.555 ;
    END
  END B[21]
  PIN B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END B[22]
  PIN B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END B[23]
  PIN B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 119.555 80.410 123.555 ;
    END
  END B[24]
  PIN B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END B[25]
  PIN B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 119.555 107.090 123.555 ;
    END
  END B[26]
  PIN B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END B[27]
  PIN B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 119.555 41.770 123.555 ;
    END
  END B[28]
  PIN B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 119.555 17.850 123.555 ;
    END
  END B[29]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 119.555 38.090 123.555 ;
    END
  END B[2]
  PIN B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 119.555 62.010 123.555 ;
    END
  END B[30]
  PIN B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END B[31]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 119.555 112.610 123.555 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 119.555 8.650 123.555 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 119.555 68.450 123.555 ;
    END
  END B[9]
  PIN Enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 100.680 112.835 101.280 ;
    END
  END Enable
  PIN Result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 119.555 95.130 123.555 ;
    END
  END Result[0]
  PIN Result[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 119.555 23.370 123.555 ;
    END
  END Result[10]
  PIN Result[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 119.555 47.290 123.555 ;
    END
  END Result[11]
  PIN Result[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 119.555 56.490 123.555 ;
    END
  END Result[12]
  PIN Result[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END Result[13]
  PIN Result[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 119.555 35.330 123.555 ;
    END
  END Result[14]
  PIN Result[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 21.800 112.835 22.400 ;
    END
  END Result[15]
  PIN Result[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END Result[16]
  PIN Result[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END Result[17]
  PIN Result[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END Result[18]
  PIN Result[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 29.960 112.835 30.560 ;
    END
  END Result[19]
  PIN Result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END Result[1]
  PIN Result[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 8.200 112.835 8.800 ;
    END
  END Result[20]
  PIN Result[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END Result[21]
  PIN Result[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END Result[22]
  PIN Result[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 53.080 112.835 53.680 ;
    END
  END Result[23]
  PIN Result[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 114.280 112.835 114.880 ;
    END
  END Result[24]
  PIN Result[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END Result[25]
  PIN Result[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 0.040 112.835 0.640 ;
    END
  END Result[26]
  PIN Result[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END Result[27]
  PIN Result[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END Result[28]
  PIN Result[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 119.555 59.250 123.555 ;
    END
  END Result[29]
  PIN Result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END Result[2]
  PIN Result[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END Result[30]
  PIN Result[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END Result[31]
  PIN Result[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END Result[32]
  PIN Result[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 78.920 112.835 79.520 ;
    END
  END Result[33]
  PIN Result[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 43.560 112.835 44.160 ;
    END
  END Result[34]
  PIN Result[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END Result[35]
  PIN Result[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END Result[36]
  PIN Result[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 12.280 112.835 12.880 ;
    END
  END Result[37]
  PIN Result[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END Result[38]
  PIN Result[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 57.160 112.835 57.760 ;
    END
  END Result[39]
  PIN Result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 96.600 112.835 97.200 ;
    END
  END Result[3]
  PIN Result[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END Result[40]
  PIN Result[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 106.120 112.835 106.720 ;
    END
  END Result[41]
  PIN Result[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 119.555 3.130 123.555 ;
    END
  END Result[42]
  PIN Result[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END Result[43]
  PIN Result[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END Result[44]
  PIN Result[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END Result[45]
  PIN Result[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END Result[46]
  PIN Result[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 119.555 11.410 123.555 ;
    END
  END Result[47]
  PIN Result[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 119.555 44.530 123.555 ;
    END
  END Result[48]
  PIN Result[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 119.555 77.650 123.555 ;
    END
  END Result[49]
  PIN Result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END Result[4]
  PIN Result[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END Result[50]
  PIN Result[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END Result[51]
  PIN Result[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 119.555 92.370 123.555 ;
    END
  END Result[52]
  PIN Result[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 119.555 71.210 123.555 ;
    END
  END Result[53]
  PIN Result[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END Result[54]
  PIN Result[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 119.555 104.330 123.555 ;
    END
  END Result[55]
  PIN Result[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 4.120 112.835 4.720 ;
    END
  END Result[56]
  PIN Result[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 119.555 5.890 123.555 ;
    END
  END Result[57]
  PIN Result[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END Result[58]
  PIN Result[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END Result[59]
  PIN Result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END Result[5]
  PIN Result[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END Result[60]
  PIN Result[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 70.760 112.835 71.360 ;
    END
  END Result[61]
  PIN Result[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END Result[62]
  PIN Result[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 119.555 89.610 123.555 ;
    END
  END Result[63]
  PIN Result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 119.555 85.930 123.555 ;
    END
  END Result[6]
  PIN Result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 119.555 14.170 123.555 ;
    END
  END Result[7]
  PIN Result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 119.555 32.570 123.555 ;
    END
  END Result[8]
  PIN Result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END Result[9]
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 43.385 107.180 44.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 76.930 107.180 78.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.605 10.640 40.205 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.490 10.640 74.090 111.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.615 107.180 28.215 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 60.160 107.180 61.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 93.705 107.180 95.305 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.665 10.640 23.265 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.550 10.640 57.150 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.435 10.640 91.035 111.760 ;
    END
  END VPWR
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.835 47.640 112.835 48.240 ;
    END
  END opcode[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.415 111.605 ;
      LAYER met1 ;
        RECT 0.070 9.900 112.630 112.500 ;
      LAYER met2 ;
        RECT 0.100 119.275 2.570 122.925 ;
        RECT 3.410 119.275 5.330 122.925 ;
        RECT 6.170 119.275 8.090 122.925 ;
        RECT 8.930 119.275 10.850 122.925 ;
        RECT 11.690 119.275 13.610 122.925 ;
        RECT 14.450 119.275 17.290 122.925 ;
        RECT 18.130 119.275 20.050 122.925 ;
        RECT 20.890 119.275 22.810 122.925 ;
        RECT 23.650 119.275 25.570 122.925 ;
        RECT 26.410 119.275 29.250 122.925 ;
        RECT 30.090 119.275 32.010 122.925 ;
        RECT 32.850 119.275 34.770 122.925 ;
        RECT 35.610 119.275 37.530 122.925 ;
        RECT 38.370 119.275 41.210 122.925 ;
        RECT 42.050 119.275 43.970 122.925 ;
        RECT 44.810 119.275 46.730 122.925 ;
        RECT 47.570 119.275 49.490 122.925 ;
        RECT 50.330 119.275 53.170 122.925 ;
        RECT 54.010 119.275 55.930 122.925 ;
        RECT 56.770 119.275 58.690 122.925 ;
        RECT 59.530 119.275 61.450 122.925 ;
        RECT 62.290 119.275 65.130 122.925 ;
        RECT 65.970 119.275 67.890 122.925 ;
        RECT 68.730 119.275 70.650 122.925 ;
        RECT 71.490 119.275 73.410 122.925 ;
        RECT 74.250 119.275 77.090 122.925 ;
        RECT 77.930 119.275 79.850 122.925 ;
        RECT 80.690 119.275 82.610 122.925 ;
        RECT 83.450 119.275 85.370 122.925 ;
        RECT 86.210 119.275 89.050 122.925 ;
        RECT 89.890 119.275 91.810 122.925 ;
        RECT 92.650 119.275 94.570 122.925 ;
        RECT 95.410 119.275 97.330 122.925 ;
        RECT 98.170 119.275 101.010 122.925 ;
        RECT 101.850 119.275 103.770 122.925 ;
        RECT 104.610 119.275 106.530 122.925 ;
        RECT 107.370 119.275 109.290 122.925 ;
        RECT 110.130 119.275 112.050 122.925 ;
        RECT 0.100 4.280 112.600 119.275 ;
        RECT 0.650 0.155 2.570 4.280 ;
        RECT 3.410 0.155 5.330 4.280 ;
        RECT 6.170 0.155 8.090 4.280 ;
        RECT 8.930 0.155 10.850 4.280 ;
        RECT 11.690 0.155 14.530 4.280 ;
        RECT 15.370 0.155 17.290 4.280 ;
        RECT 18.130 0.155 20.050 4.280 ;
        RECT 20.890 0.155 22.810 4.280 ;
        RECT 23.650 0.155 26.490 4.280 ;
        RECT 27.330 0.155 29.250 4.280 ;
        RECT 30.090 0.155 32.010 4.280 ;
        RECT 32.850 0.155 34.770 4.280 ;
        RECT 35.610 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.210 4.280 ;
        RECT 42.050 0.155 43.970 4.280 ;
        RECT 44.810 0.155 46.730 4.280 ;
        RECT 47.570 0.155 50.410 4.280 ;
        RECT 51.250 0.155 53.170 4.280 ;
        RECT 54.010 0.155 55.930 4.280 ;
        RECT 56.770 0.155 58.690 4.280 ;
        RECT 59.530 0.155 62.370 4.280 ;
        RECT 63.210 0.155 65.130 4.280 ;
        RECT 65.970 0.155 67.890 4.280 ;
        RECT 68.730 0.155 70.650 4.280 ;
        RECT 71.490 0.155 74.330 4.280 ;
        RECT 75.170 0.155 77.090 4.280 ;
        RECT 77.930 0.155 79.850 4.280 ;
        RECT 80.690 0.155 82.610 4.280 ;
        RECT 83.450 0.155 86.290 4.280 ;
        RECT 87.130 0.155 89.050 4.280 ;
        RECT 89.890 0.155 91.810 4.280 ;
        RECT 92.650 0.155 94.570 4.280 ;
        RECT 95.410 0.155 98.250 4.280 ;
        RECT 99.090 0.155 101.010 4.280 ;
        RECT 101.850 0.155 103.770 4.280 ;
        RECT 104.610 0.155 106.530 4.280 ;
        RECT 107.370 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 122.040 108.835 122.905 ;
        RECT 4.000 119.360 108.835 122.040 ;
        RECT 4.400 117.960 108.435 119.360 ;
        RECT 4.000 115.280 108.835 117.960 ;
        RECT 4.400 113.880 108.435 115.280 ;
        RECT 4.000 111.200 108.835 113.880 ;
        RECT 4.400 109.800 108.435 111.200 ;
        RECT 4.000 107.120 108.835 109.800 ;
        RECT 4.000 105.760 108.435 107.120 ;
        RECT 4.400 105.720 108.435 105.760 ;
        RECT 4.400 104.360 108.835 105.720 ;
        RECT 4.000 101.680 108.835 104.360 ;
        RECT 4.400 100.280 108.435 101.680 ;
        RECT 4.000 97.600 108.835 100.280 ;
        RECT 4.400 96.200 108.435 97.600 ;
        RECT 4.000 93.520 108.835 96.200 ;
        RECT 4.400 92.120 108.435 93.520 ;
        RECT 4.000 89.440 108.835 92.120 ;
        RECT 4.000 88.080 108.435 89.440 ;
        RECT 4.400 88.040 108.435 88.080 ;
        RECT 4.400 86.680 108.835 88.040 ;
        RECT 4.000 84.000 108.835 86.680 ;
        RECT 4.400 82.600 108.435 84.000 ;
        RECT 4.000 79.920 108.835 82.600 ;
        RECT 4.400 78.520 108.435 79.920 ;
        RECT 4.000 75.840 108.835 78.520 ;
        RECT 4.400 74.440 108.435 75.840 ;
        RECT 4.000 71.760 108.835 74.440 ;
        RECT 4.000 70.400 108.435 71.760 ;
        RECT 4.400 70.360 108.435 70.400 ;
        RECT 4.400 69.000 108.835 70.360 ;
        RECT 4.000 66.320 108.835 69.000 ;
        RECT 4.400 64.920 108.435 66.320 ;
        RECT 4.000 62.240 108.835 64.920 ;
        RECT 4.400 60.840 108.435 62.240 ;
        RECT 4.000 58.160 108.835 60.840 ;
        RECT 4.400 56.760 108.435 58.160 ;
        RECT 4.000 54.080 108.835 56.760 ;
        RECT 4.000 52.720 108.435 54.080 ;
        RECT 4.400 52.680 108.435 52.720 ;
        RECT 4.400 51.320 108.835 52.680 ;
        RECT 4.000 48.640 108.835 51.320 ;
        RECT 4.400 47.240 108.435 48.640 ;
        RECT 4.000 44.560 108.835 47.240 ;
        RECT 4.400 43.160 108.435 44.560 ;
        RECT 4.000 40.480 108.835 43.160 ;
        RECT 4.400 39.080 108.435 40.480 ;
        RECT 4.000 36.400 108.835 39.080 ;
        RECT 4.000 35.040 108.435 36.400 ;
        RECT 4.400 35.000 108.435 35.040 ;
        RECT 4.400 33.640 108.835 35.000 ;
        RECT 4.000 30.960 108.835 33.640 ;
        RECT 4.400 29.560 108.435 30.960 ;
        RECT 4.000 26.880 108.835 29.560 ;
        RECT 4.400 25.480 108.435 26.880 ;
        RECT 4.000 22.800 108.835 25.480 ;
        RECT 4.400 21.400 108.435 22.800 ;
        RECT 4.000 18.720 108.835 21.400 ;
        RECT 4.000 17.360 108.435 18.720 ;
        RECT 4.400 17.320 108.435 17.360 ;
        RECT 4.400 15.960 108.835 17.320 ;
        RECT 4.000 13.280 108.835 15.960 ;
        RECT 4.400 11.880 108.435 13.280 ;
        RECT 4.000 9.200 108.835 11.880 ;
        RECT 4.400 7.800 108.435 9.200 ;
        RECT 4.000 5.120 108.835 7.800 ;
        RECT 4.400 3.720 108.435 5.120 ;
        RECT 4.000 1.040 108.835 3.720 ;
        RECT 4.000 0.175 108.435 1.040 ;
      LAYER met4 ;
        RECT 23.665 10.640 38.205 111.760 ;
        RECT 40.605 10.640 55.150 111.760 ;
        RECT 57.550 10.640 72.090 111.760 ;
        RECT 74.490 10.640 89.035 111.760 ;
        RECT 91.435 10.640 102.745 111.760 ;
  END
END alu32
END LIBRARY

